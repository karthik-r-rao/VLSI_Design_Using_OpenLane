magic
tech sky130A
magscale 1 2
timestamp 1618160920
<< obsli1 >>
rect 1104 1785 85192 85969
<< obsm1 >>
rect 1104 1572 85192 86148
<< metal2 >>
rect 1398 87660 1454 88460
rect 3238 87660 3294 88460
rect 5078 87660 5134 88460
rect 6918 87660 6974 88460
rect 8298 87660 8354 88460
rect 10138 87660 10194 88460
rect 11978 87660 12034 88460
rect 13358 87660 13414 88460
rect 15198 87660 15254 88460
rect 17038 87660 17094 88460
rect 18878 87660 18934 88460
rect 20258 87660 20314 88460
rect 22098 87660 22154 88460
rect 23938 87660 23994 88460
rect 25778 87660 25834 88460
rect 27158 87660 27214 88460
rect 28998 87660 29054 88460
rect 30838 87660 30894 88460
rect 32678 87660 32734 88460
rect 34058 87660 34114 88460
rect 35898 87660 35954 88460
rect 37738 87660 37794 88460
rect 39578 87660 39634 88460
rect 40958 87660 41014 88460
rect 42798 87660 42854 88460
rect 44638 87660 44694 88460
rect 46478 87660 46534 88460
rect 47858 87660 47914 88460
rect 49698 87660 49754 88460
rect 51538 87660 51594 88460
rect 52918 87660 52974 88460
rect 54758 87660 54814 88460
rect 56598 87660 56654 88460
rect 58438 87660 58494 88460
rect 59818 87660 59874 88460
rect 61658 87660 61714 88460
rect 63498 87660 63554 88460
rect 65338 87660 65394 88460
rect 66718 87660 66774 88460
rect 68558 87660 68614 88460
rect 70398 87660 70454 88460
rect 72238 87660 72294 88460
rect 73618 87660 73674 88460
rect 75458 87660 75514 88460
rect 77298 87660 77354 88460
rect 79138 87660 79194 88460
rect 80518 87660 80574 88460
rect 82358 87660 82414 88460
rect 84198 87660 84254 88460
rect 85578 87660 85634 88460
rect 478 0 534 800
rect 1858 0 1914 800
rect 3698 0 3754 800
rect 5538 0 5594 800
rect 6918 0 6974 800
rect 8758 0 8814 800
rect 10598 0 10654 800
rect 12438 0 12494 800
rect 13818 0 13874 800
rect 15658 0 15714 800
rect 17498 0 17554 800
rect 19338 0 19394 800
rect 20718 0 20774 800
rect 22558 0 22614 800
rect 24398 0 24454 800
rect 26238 0 26294 800
rect 27618 0 27674 800
rect 29458 0 29514 800
rect 31298 0 31354 800
rect 33138 0 33194 800
rect 34518 0 34574 800
rect 36358 0 36414 800
rect 38198 0 38254 800
rect 39578 0 39634 800
rect 41418 0 41474 800
rect 43258 0 43314 800
rect 45098 0 45154 800
rect 46478 0 46534 800
rect 48318 0 48374 800
rect 50158 0 50214 800
rect 51998 0 52054 800
rect 53378 0 53434 800
rect 55218 0 55274 800
rect 57058 0 57114 800
rect 58898 0 58954 800
rect 60278 0 60334 800
rect 62118 0 62174 800
rect 63958 0 64014 800
rect 65798 0 65854 800
rect 67178 0 67234 800
rect 69018 0 69074 800
rect 70858 0 70914 800
rect 72698 0 72754 800
rect 74078 0 74134 800
rect 75918 0 75974 800
rect 77758 0 77814 800
rect 79138 0 79194 800
rect 80978 0 81034 800
rect 82818 0 82874 800
rect 84658 0 84714 800
<< obsm2 >>
rect 478 87604 1342 87660
rect 1510 87604 3182 87660
rect 3350 87604 5022 87660
rect 5190 87604 6862 87660
rect 7030 87604 8242 87660
rect 8410 87604 10082 87660
rect 10250 87604 11922 87660
rect 12090 87604 13302 87660
rect 13470 87604 15142 87660
rect 15310 87604 16982 87660
rect 17150 87604 18822 87660
rect 18990 87604 20202 87660
rect 20370 87604 22042 87660
rect 22210 87604 23882 87660
rect 24050 87604 25722 87660
rect 25890 87604 27102 87660
rect 27270 87604 28942 87660
rect 29110 87604 30782 87660
rect 30950 87604 32622 87660
rect 32790 87604 34002 87660
rect 34170 87604 35842 87660
rect 36010 87604 37682 87660
rect 37850 87604 39522 87660
rect 39690 87604 40902 87660
rect 41070 87604 42742 87660
rect 42910 87604 44582 87660
rect 44750 87604 46422 87660
rect 46590 87604 47802 87660
rect 47970 87604 49642 87660
rect 49810 87604 51482 87660
rect 51650 87604 52862 87660
rect 53030 87604 54702 87660
rect 54870 87604 56542 87660
rect 56710 87604 58382 87660
rect 58550 87604 59762 87660
rect 59930 87604 61602 87660
rect 61770 87604 63442 87660
rect 63610 87604 65282 87660
rect 65450 87604 66662 87660
rect 66830 87604 68502 87660
rect 68670 87604 70342 87660
rect 70510 87604 72182 87660
rect 72350 87604 73562 87660
rect 73730 87604 75402 87660
rect 75570 87604 77242 87660
rect 77410 87604 79082 87660
rect 79250 87604 80462 87660
rect 80630 87604 82302 87660
rect 82470 87604 84142 87660
rect 84310 87604 85522 87660
rect 478 856 85620 87604
rect 590 711 1802 856
rect 1970 711 3642 856
rect 3810 711 5482 856
rect 5650 711 6862 856
rect 7030 711 8702 856
rect 8870 711 10542 856
rect 10710 711 12382 856
rect 12550 711 13762 856
rect 13930 711 15602 856
rect 15770 711 17442 856
rect 17610 711 19282 856
rect 19450 711 20662 856
rect 20830 711 22502 856
rect 22670 711 24342 856
rect 24510 711 26182 856
rect 26350 711 27562 856
rect 27730 711 29402 856
rect 29570 711 31242 856
rect 31410 711 33082 856
rect 33250 711 34462 856
rect 34630 711 36302 856
rect 36470 711 38142 856
rect 38310 711 39522 856
rect 39690 711 41362 856
rect 41530 711 43202 856
rect 43370 711 45042 856
rect 45210 711 46422 856
rect 46590 711 48262 856
rect 48430 711 50102 856
rect 50270 711 51942 856
rect 52110 711 53322 856
rect 53490 711 55162 856
rect 55330 711 57002 856
rect 57170 711 58842 856
rect 59010 711 60222 856
rect 60390 711 62062 856
rect 62230 711 63902 856
rect 64070 711 65742 856
rect 65910 711 67122 856
rect 67290 711 68962 856
rect 69130 711 70802 856
rect 70970 711 72642 856
rect 72810 711 74022 856
rect 74190 711 75862 856
rect 76030 711 77702 856
rect 77870 711 79082 856
rect 79250 711 80922 856
rect 81090 711 82762 856
rect 82930 711 84602 856
rect 84770 711 85620 856
<< metal3 >>
rect 0 87048 800 87168
rect 85516 85008 86316 85128
rect 0 84328 800 84448
rect 85516 82288 86316 82408
rect 0 81608 800 81728
rect 85516 79568 86316 79688
rect 0 78888 800 79008
rect 85516 77528 86316 77648
rect 0 76848 800 76968
rect 85516 74808 86316 74928
rect 0 74128 800 74248
rect 85516 72088 86316 72208
rect 0 71408 800 71528
rect 85516 69368 86316 69488
rect 0 68688 800 68808
rect 85516 67328 86316 67448
rect 0 66648 800 66768
rect 85516 64608 86316 64728
rect 0 63928 800 64048
rect 85516 61888 86316 62008
rect 0 61208 800 61328
rect 85516 59168 86316 59288
rect 0 58488 800 58608
rect 85516 57128 86316 57248
rect 0 56448 800 56568
rect 85516 54408 86316 54528
rect 0 53728 800 53848
rect 85516 51688 86316 51808
rect 0 51008 800 51128
rect 0 48968 800 49088
rect 85516 48968 86316 49088
rect 85516 46928 86316 47048
rect 0 46248 800 46368
rect 85516 44208 86316 44328
rect 0 43528 800 43648
rect 85516 41488 86316 41608
rect 0 40808 800 40928
rect 0 38768 800 38888
rect 85516 38768 86316 38888
rect 85516 36728 86316 36848
rect 0 36048 800 36168
rect 85516 34008 86316 34128
rect 0 33328 800 33448
rect 85516 31288 86316 31408
rect 0 30608 800 30728
rect 85516 29248 86316 29368
rect 0 28568 800 28688
rect 85516 26528 86316 26648
rect 0 25848 800 25968
rect 85516 23808 86316 23928
rect 0 23128 800 23248
rect 85516 21088 86316 21208
rect 0 20408 800 20528
rect 85516 19048 86316 19168
rect 0 18368 800 18488
rect 85516 16328 86316 16448
rect 0 15648 800 15768
rect 85516 13608 86316 13728
rect 0 12928 800 13048
rect 85516 10888 86316 11008
rect 0 10208 800 10328
rect 85516 8848 86316 8968
rect 0 8168 800 8288
rect 85516 6128 86316 6248
rect 0 5448 800 5568
rect 85516 3408 86316 3528
rect 0 2728 800 2848
rect 85516 688 86316 808
<< obsm3 >>
rect 880 86968 85516 87141
rect 473 85208 85516 86968
rect 473 84928 85436 85208
rect 473 84528 85516 84928
rect 880 84248 85516 84528
rect 473 82488 85516 84248
rect 473 82208 85436 82488
rect 473 81808 85516 82208
rect 880 81528 85516 81808
rect 473 79768 85516 81528
rect 473 79488 85436 79768
rect 473 79088 85516 79488
rect 880 78808 85516 79088
rect 473 77728 85516 78808
rect 473 77448 85436 77728
rect 473 77048 85516 77448
rect 880 76768 85516 77048
rect 473 75008 85516 76768
rect 473 74728 85436 75008
rect 473 74328 85516 74728
rect 880 74048 85516 74328
rect 473 72288 85516 74048
rect 473 72008 85436 72288
rect 473 71608 85516 72008
rect 880 71328 85516 71608
rect 473 69568 85516 71328
rect 473 69288 85436 69568
rect 473 68888 85516 69288
rect 880 68608 85516 68888
rect 473 67528 85516 68608
rect 473 67248 85436 67528
rect 473 66848 85516 67248
rect 880 66568 85516 66848
rect 473 64808 85516 66568
rect 473 64528 85436 64808
rect 473 64128 85516 64528
rect 880 63848 85516 64128
rect 473 62088 85516 63848
rect 473 61808 85436 62088
rect 473 61408 85516 61808
rect 880 61128 85516 61408
rect 473 59368 85516 61128
rect 473 59088 85436 59368
rect 473 58688 85516 59088
rect 880 58408 85516 58688
rect 473 57328 85516 58408
rect 473 57048 85436 57328
rect 473 56648 85516 57048
rect 880 56368 85516 56648
rect 473 54608 85516 56368
rect 473 54328 85436 54608
rect 473 53928 85516 54328
rect 880 53648 85516 53928
rect 473 51888 85516 53648
rect 473 51608 85436 51888
rect 473 51208 85516 51608
rect 880 50928 85516 51208
rect 473 49168 85516 50928
rect 880 48888 85436 49168
rect 473 47128 85516 48888
rect 473 46848 85436 47128
rect 473 46448 85516 46848
rect 880 46168 85516 46448
rect 473 44408 85516 46168
rect 473 44128 85436 44408
rect 473 43728 85516 44128
rect 880 43448 85516 43728
rect 473 41688 85516 43448
rect 473 41408 85436 41688
rect 473 41008 85516 41408
rect 880 40728 85516 41008
rect 473 38968 85516 40728
rect 880 38688 85436 38968
rect 473 36928 85516 38688
rect 473 36648 85436 36928
rect 473 36248 85516 36648
rect 880 35968 85516 36248
rect 473 34208 85516 35968
rect 473 33928 85436 34208
rect 473 33528 85516 33928
rect 880 33248 85516 33528
rect 473 31488 85516 33248
rect 473 31208 85436 31488
rect 473 30808 85516 31208
rect 880 30528 85516 30808
rect 473 29448 85516 30528
rect 473 29168 85436 29448
rect 473 28768 85516 29168
rect 880 28488 85516 28768
rect 473 26728 85516 28488
rect 473 26448 85436 26728
rect 473 26048 85516 26448
rect 880 25768 85516 26048
rect 473 24008 85516 25768
rect 473 23728 85436 24008
rect 473 23328 85516 23728
rect 880 23048 85516 23328
rect 473 21288 85516 23048
rect 473 21008 85436 21288
rect 473 20608 85516 21008
rect 880 20328 85516 20608
rect 473 19248 85516 20328
rect 473 18968 85436 19248
rect 473 18568 85516 18968
rect 880 18288 85516 18568
rect 473 16528 85516 18288
rect 473 16248 85436 16528
rect 473 15848 85516 16248
rect 880 15568 85516 15848
rect 473 13808 85516 15568
rect 473 13528 85436 13808
rect 473 13128 85516 13528
rect 880 12848 85516 13128
rect 473 11088 85516 12848
rect 473 10808 85436 11088
rect 473 10408 85516 10808
rect 880 10128 85516 10408
rect 473 9048 85516 10128
rect 473 8768 85436 9048
rect 473 8368 85516 8768
rect 880 8088 85516 8368
rect 473 6328 85516 8088
rect 473 6048 85436 6328
rect 473 5648 85516 6048
rect 880 5368 85516 5648
rect 473 3608 85516 5368
rect 473 3328 85436 3608
rect 473 2928 85516 3328
rect 880 2648 85516 2928
rect 473 888 85516 2648
rect 473 715 85436 888
<< metal4 >>
rect 4208 2128 4528 86000
rect 19568 2128 19888 86000
rect 34928 2128 35248 86000
rect 50288 2128 50608 86000
rect 65648 2128 65968 86000
rect 81008 2128 81328 86000
<< obsm4 >>
rect 1814 2619 4128 85645
rect 4608 2619 19488 85645
rect 19968 2619 34848 85645
rect 35328 2619 50208 85645
rect 50688 2619 65568 85645
rect 66048 2619 80928 85645
rect 81408 2619 82557 85645
<< metal5 >>
rect 1104 81888 85192 82208
rect 1104 66570 85192 66890
rect 1104 51252 85192 51572
rect 1104 35934 85192 36254
rect 1104 20616 85192 20936
rect 1104 5298 85192 5618
<< obsm5 >>
rect 1772 36574 78636 48100
rect 1772 21256 78636 35614
rect 1772 5938 78636 20296
rect 1772 3580 78636 4978
<< labels >>
rlabel metal2 s 77298 87660 77354 88460 6 clk
port 1 nsew signal input
rlabel metal2 s 6918 87660 6974 88460 6 data_address[0]
port 2 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 data_address[10]
port 3 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 data_address[11]
port 4 nsew signal output
rlabel metal2 s 82358 87660 82414 88460 6 data_address[12]
port 5 nsew signal output
rlabel metal2 s 30838 87660 30894 88460 6 data_address[13]
port 6 nsew signal output
rlabel metal2 s 70398 87660 70454 88460 6 data_address[14]
port 7 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 data_address[15]
port 8 nsew signal output
rlabel metal2 s 10138 87660 10194 88460 6 data_address[16]
port 9 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 data_address[17]
port 10 nsew signal output
rlabel metal2 s 66718 87660 66774 88460 6 data_address[18]
port 11 nsew signal output
rlabel metal2 s 85578 87660 85634 88460 6 data_address[19]
port 12 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 data_address[1]
port 13 nsew signal output
rlabel metal3 s 85516 8848 86316 8968 6 data_address[20]
port 14 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 data_address[21]
port 15 nsew signal output
rlabel metal2 s 39578 87660 39634 88460 6 data_address[22]
port 16 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 data_address[23]
port 17 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 data_address[24]
port 18 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 data_address[25]
port 19 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 data_address[26]
port 20 nsew signal output
rlabel metal2 s 51538 87660 51594 88460 6 data_address[27]
port 21 nsew signal output
rlabel metal2 s 17038 87660 17094 88460 6 data_address[28]
port 22 nsew signal output
rlabel metal2 s 68558 87660 68614 88460 6 data_address[29]
port 23 nsew signal output
rlabel metal2 s 63498 87660 63554 88460 6 data_address[2]
port 24 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 data_address[30]
port 25 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 data_address[31]
port 26 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 data_address[3]
port 27 nsew signal output
rlabel metal2 s 1398 87660 1454 88460 6 data_address[4]
port 28 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 data_address[5]
port 29 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 data_address[6]
port 30 nsew signal output
rlabel metal2 s 56598 87660 56654 88460 6 data_address[7]
port 31 nsew signal output
rlabel metal3 s 85516 57128 86316 57248 6 data_address[8]
port 32 nsew signal output
rlabel metal3 s 85516 23808 86316 23928 6 data_address[9]
port 33 nsew signal output
rlabel metal3 s 85516 82288 86316 82408 6 instruction[0]
port 34 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 instruction[10]
port 35 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 instruction[11]
port 36 nsew signal input
rlabel metal3 s 85516 74808 86316 74928 6 instruction[12]
port 37 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 instruction[13]
port 38 nsew signal input
rlabel metal3 s 85516 31288 86316 31408 6 instruction[14]
port 39 nsew signal input
rlabel metal2 s 15198 87660 15254 88460 6 instruction[15]
port 40 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 instruction[16]
port 41 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 instruction[17]
port 42 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 instruction[18]
port 43 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 instruction[19]
port 44 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 instruction[1]
port 45 nsew signal input
rlabel metal3 s 85516 79568 86316 79688 6 instruction[20]
port 46 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 instruction[21]
port 47 nsew signal input
rlabel metal3 s 85516 688 86316 808 6 instruction[22]
port 48 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 instruction[23]
port 49 nsew signal input
rlabel metal3 s 85516 77528 86316 77648 6 instruction[24]
port 50 nsew signal input
rlabel metal2 s 8298 87660 8354 88460 6 instruction[25]
port 51 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 instruction[26]
port 52 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 instruction[27]
port 53 nsew signal input
rlabel metal2 s 34058 87660 34114 88460 6 instruction[28]
port 54 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 instruction[29]
port 55 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 instruction[2]
port 56 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 instruction[30]
port 57 nsew signal input
rlabel metal2 s 13358 87660 13414 88460 6 instruction[31]
port 58 nsew signal input
rlabel metal3 s 85516 21088 86316 21208 6 instruction[3]
port 59 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 instruction[4]
port 60 nsew signal input
rlabel metal3 s 85516 6128 86316 6248 6 instruction[5]
port 61 nsew signal input
rlabel metal3 s 85516 26528 86316 26648 6 instruction[6]
port 62 nsew signal input
rlabel metal2 s 22098 87660 22154 88460 6 instruction[7]
port 63 nsew signal input
rlabel metal2 s 54758 87660 54814 88460 6 instruction[8]
port 64 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 instruction[9]
port 65 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 pc[0]
port 66 nsew signal output
rlabel metal2 s 37738 87660 37794 88460 6 pc[10]
port 67 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 pc[11]
port 68 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 pc[12]
port 69 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 pc[13]
port 70 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 pc[14]
port 71 nsew signal output
rlabel metal3 s 85516 46928 86316 47048 6 pc[15]
port 72 nsew signal output
rlabel metal2 s 52918 87660 52974 88460 6 pc[16]
port 73 nsew signal output
rlabel metal2 s 23938 87660 23994 88460 6 pc[17]
port 74 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 pc[18]
port 75 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 pc[19]
port 76 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 pc[1]
port 77 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 pc[20]
port 78 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 pc[21]
port 79 nsew signal output
rlabel metal2 s 58438 87660 58494 88460 6 pc[22]
port 80 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 pc[23]
port 81 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 pc[24]
port 82 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 pc[25]
port 83 nsew signal output
rlabel metal2 s 20258 87660 20314 88460 6 pc[26]
port 84 nsew signal output
rlabel metal2 s 18878 87660 18934 88460 6 pc[27]
port 85 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 pc[28]
port 86 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 pc[29]
port 87 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 pc[2]
port 88 nsew signal output
rlabel metal2 s 75458 87660 75514 88460 6 pc[30]
port 89 nsew signal output
rlabel metal3 s 85516 51688 86316 51808 6 pc[31]
port 90 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 pc[3]
port 91 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 pc[4]
port 92 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 pc[5]
port 93 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 pc[6]
port 94 nsew signal output
rlabel metal3 s 85516 67328 86316 67448 6 pc[7]
port 95 nsew signal output
rlabel metal3 s 85516 16328 86316 16448 6 pc[8]
port 96 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 pc[9]
port 97 nsew signal output
rlabel metal2 s 5078 87660 5134 88460 6 rdata[0]
port 98 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 rdata[10]
port 99 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 rdata[11]
port 100 nsew signal input
rlabel metal3 s 85516 54408 86316 54528 6 rdata[12]
port 101 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 rdata[13]
port 102 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 rdata[14]
port 103 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 rdata[15]
port 104 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 rdata[16]
port 105 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 rdata[17]
port 106 nsew signal input
rlabel metal3 s 85516 41488 86316 41608 6 rdata[18]
port 107 nsew signal input
rlabel metal2 s 35898 87660 35954 88460 6 rdata[19]
port 108 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 rdata[1]
port 109 nsew signal input
rlabel metal2 s 40958 87660 41014 88460 6 rdata[20]
port 110 nsew signal input
rlabel metal2 s 80518 87660 80574 88460 6 rdata[21]
port 111 nsew signal input
rlabel metal3 s 85516 85008 86316 85128 6 rdata[22]
port 112 nsew signal input
rlabel metal3 s 85516 44208 86316 44328 6 rdata[23]
port 113 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 rdata[24]
port 114 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 rdata[25]
port 115 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 rdata[26]
port 116 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 rdata[27]
port 117 nsew signal input
rlabel metal3 s 85516 38768 86316 38888 6 rdata[28]
port 118 nsew signal input
rlabel metal2 s 49698 87660 49754 88460 6 rdata[29]
port 119 nsew signal input
rlabel metal3 s 85516 59168 86316 59288 6 rdata[2]
port 120 nsew signal input
rlabel metal2 s 84198 87660 84254 88460 6 rdata[30]
port 121 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 rdata[31]
port 122 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 rdata[3]
port 123 nsew signal input
rlabel metal3 s 85516 29248 86316 29368 6 rdata[4]
port 124 nsew signal input
rlabel metal3 s 85516 19048 86316 19168 6 rdata[5]
port 125 nsew signal input
rlabel metal2 s 25778 87660 25834 88460 6 rdata[6]
port 126 nsew signal input
rlabel metal2 s 3238 87660 3294 88460 6 rdata[7]
port 127 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 rdata[8]
port 128 nsew signal input
rlabel metal2 s 61658 87660 61714 88460 6 rdata[9]
port 129 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 ren
port 130 nsew signal output
rlabel metal3 s 85516 61888 86316 62008 6 rst
port 131 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 wdata[0]
port 132 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 wdata[10]
port 133 nsew signal output
rlabel metal2 s 11978 87660 12034 88460 6 wdata[11]
port 134 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 wdata[12]
port 135 nsew signal output
rlabel metal2 s 79138 87660 79194 88460 6 wdata[13]
port 136 nsew signal output
rlabel metal3 s 85516 34008 86316 34128 6 wdata[14]
port 137 nsew signal output
rlabel metal2 s 47858 87660 47914 88460 6 wdata[15]
port 138 nsew signal output
rlabel metal2 s 32678 87660 32734 88460 6 wdata[16]
port 139 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 wdata[17]
port 140 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wdata[18]
port 141 nsew signal output
rlabel metal3 s 85516 72088 86316 72208 6 wdata[19]
port 142 nsew signal output
rlabel metal3 s 85516 64608 86316 64728 6 wdata[1]
port 143 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wdata[20]
port 144 nsew signal output
rlabel metal2 s 65338 87660 65394 88460 6 wdata[21]
port 145 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wdata[22]
port 146 nsew signal output
rlabel metal3 s 85516 13608 86316 13728 6 wdata[23]
port 147 nsew signal output
rlabel metal2 s 28998 87660 29054 88460 6 wdata[24]
port 148 nsew signal output
rlabel metal3 s 85516 48968 86316 49088 6 wdata[25]
port 149 nsew signal output
rlabel metal3 s 85516 69368 86316 69488 6 wdata[26]
port 150 nsew signal output
rlabel metal2 s 72238 87660 72294 88460 6 wdata[27]
port 151 nsew signal output
rlabel metal2 s 59818 87660 59874 88460 6 wdata[28]
port 152 nsew signal output
rlabel metal2 s 478 0 534 800 6 wdata[29]
port 153 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wdata[2]
port 154 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 wdata[30]
port 155 nsew signal output
rlabel metal2 s 44638 87660 44694 88460 6 wdata[31]
port 156 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wdata[3]
port 157 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 wdata[4]
port 158 nsew signal output
rlabel metal2 s 73618 87660 73674 88460 6 wdata[5]
port 159 nsew signal output
rlabel metal2 s 27158 87660 27214 88460 6 wdata[6]
port 160 nsew signal output
rlabel metal3 s 85516 36728 86316 36848 6 wdata[7]
port 161 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 wdata[8]
port 162 nsew signal output
rlabel metal2 s 46478 87660 46534 88460 6 wdata[9]
port 163 nsew signal output
rlabel metal3 s 85516 10888 86316 11008 6 wen
port 164 nsew signal output
rlabel metal3 s 85516 3408 86316 3528 6 wstrobe[0]
port 165 nsew signal output
rlabel metal2 s 42798 87660 42854 88460 6 wstrobe[1]
port 166 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 wstrobe[2]
port 167 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 wstrobe[3]
port 168 nsew signal output
rlabel metal4 s 65648 2128 65968 86000 6 VPWR
port 169 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 86000 6 VPWR
port 170 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 86000 6 VPWR
port 171 nsew power bidirectional
rlabel metal5 s 1104 66570 85192 66890 6 VPWR
port 172 nsew power bidirectional
rlabel metal5 s 1104 35934 85192 36254 6 VPWR
port 173 nsew power bidirectional
rlabel metal5 s 1104 5298 85192 5618 6 VPWR
port 174 nsew power bidirectional
rlabel metal4 s 81008 2128 81328 86000 6 VGND
port 175 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 86000 6 VGND
port 176 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 86000 6 VGND
port 177 nsew ground bidirectional
rlabel metal5 s 1104 81888 85192 82208 6 VGND
port 178 nsew ground bidirectional
rlabel metal5 s 1104 51252 85192 51572 6 VGND
port 179 nsew ground bidirectional
rlabel metal5 s 1104 20616 85192 20936 6 VGND
port 180 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 86316 88460
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/core/runs/core/results/magic/core.gds
string GDS_END 26704532
string GDS_START 817428
<< end >>

