localparam LUI = 7'b0110111;
localparam AUIPC = 7'b0010111;
localparam JAL = 7'b1101111;
localparam JALR = 7'b1100111;
localparam BRANCH = 7'b1100011;
localparam LOAD = 7'b0000011;
localparam STORE = 7'b0100011;
localparam IMM = 7'b0010011;
localparam REG = 7'b0110011;

localparam BEQ = 3'b000; 
localparam BNE = 3'b001;
localparam BLT = 3'b100;
localparam BGE = 3'b101;
localparam BLTU = 3'b110;
localparam BGEU = 3'b111;
localparam LB = 3'b000;
localparam LH = 3'b001;
localparam LW = 3'b010;
localparam LBU = 3'b100;
localparam LHU = 3'b101;
localparam SB = 3'b000;
localparam SH = 3'b001;
localparam SW = 3'b010;
localparam ADDI = 3'b000;
localparam SLTI = 3'b010;
localparam SLTIU = 3'b011;
localparam XORI = 3'b100;
localparam ORI = 3'b110;
localparam ANDI = 3'b111;
localparam SLLI = 3'b001;
localparam SRI = 3'b101;    // SRLI and SRAI
localparam ADDSUB = 3'b000; // ADD and SUB  
localparam SLL = 3'b001;
localparam SLT = 3'b010;
localparam SLTU = 3'b011;
localparam XOR = 3'b100;
localparam SR = 3'b101;     // SRL and SRA
localparam OR = 3'b110;
localparam AND = 3'b111;

localparam SRLI = 7'b0000000;
localparam SRAI = 7'b0100000;
localparam ADD = 7'b0000000;
localparam SUB = 7'b0100000;
localparam SRL = 7'b0000000;
localparam SRA = 7'b0100000;