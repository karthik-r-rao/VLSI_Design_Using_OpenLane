VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 431.580 BY 442.300 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 438.300 386.770 442.300 ;
    END
  END clk
  PIN data_address[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 438.300 34.870 442.300 ;
    END
  END data_address[0]
  PIN data_address[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END data_address[10]
  PIN data_address[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END data_address[11]
  PIN data_address[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 438.300 412.070 442.300 ;
    END
  END data_address[12]
  PIN data_address[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 438.300 154.470 442.300 ;
    END
  END data_address[13]
  PIN data_address[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 438.300 352.270 442.300 ;
    END
  END data_address[14]
  PIN data_address[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END data_address[15]
  PIN data_address[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 438.300 50.970 442.300 ;
    END
  END data_address[16]
  PIN data_address[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END data_address[17]
  PIN data_address[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 438.300 333.870 442.300 ;
    END
  END data_address[18]
  PIN data_address[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 438.300 428.170 442.300 ;
    END
  END data_address[19]
  PIN data_address[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END data_address[1]
  PIN data_address[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 44.240 431.580 44.840 ;
    END
  END data_address[20]
  PIN data_address[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END data_address[21]
  PIN data_address[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 438.300 198.170 442.300 ;
    END
  END data_address[22]
  PIN data_address[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END data_address[23]
  PIN data_address[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END data_address[24]
  PIN data_address[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END data_address[25]
  PIN data_address[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END data_address[26]
  PIN data_address[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 438.300 257.970 442.300 ;
    END
  END data_address[27]
  PIN data_address[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 438.300 85.470 442.300 ;
    END
  END data_address[28]
  PIN data_address[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 438.300 343.070 442.300 ;
    END
  END data_address[29]
  PIN data_address[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 438.300 317.770 442.300 ;
    END
  END data_address[2]
  PIN data_address[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END data_address[30]
  PIN data_address[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END data_address[31]
  PIN data_address[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END data_address[3]
  PIN data_address[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 438.300 7.270 442.300 ;
    END
  END data_address[4]
  PIN data_address[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END data_address[5]
  PIN data_address[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END data_address[6]
  PIN data_address[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 438.300 283.270 442.300 ;
    END
  END data_address[7]
  PIN data_address[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 285.640 431.580 286.240 ;
    END
  END data_address[8]
  PIN data_address[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 119.040 431.580 119.640 ;
    END
  END data_address[9]
  PIN instruction[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 411.440 431.580 412.040 ;
    END
  END instruction[0]
  PIN instruction[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END instruction[10]
  PIN instruction[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END instruction[11]
  PIN instruction[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 374.040 431.580 374.640 ;
    END
  END instruction[12]
  PIN instruction[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END instruction[13]
  PIN instruction[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 156.440 431.580 157.040 ;
    END
  END instruction[14]
  PIN instruction[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 438.300 76.270 442.300 ;
    END
  END instruction[15]
  PIN instruction[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END instruction[16]
  PIN instruction[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END instruction[17]
  PIN instruction[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END instruction[18]
  PIN instruction[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END instruction[19]
  PIN instruction[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END instruction[1]
  PIN instruction[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 397.840 431.580 398.440 ;
    END
  END instruction[20]
  PIN instruction[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END instruction[21]
  PIN instruction[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 3.440 431.580 4.040 ;
    END
  END instruction[22]
  PIN instruction[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END instruction[23]
  PIN instruction[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 387.640 431.580 388.240 ;
    END
  END instruction[24]
  PIN instruction[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 438.300 41.770 442.300 ;
    END
  END instruction[25]
  PIN instruction[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END instruction[26]
  PIN instruction[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END instruction[27]
  PIN instruction[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 438.300 170.570 442.300 ;
    END
  END instruction[28]
  PIN instruction[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END instruction[29]
  PIN instruction[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END instruction[2]
  PIN instruction[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END instruction[30]
  PIN instruction[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 438.300 67.070 442.300 ;
    END
  END instruction[31]
  PIN instruction[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 105.440 431.580 106.040 ;
    END
  END instruction[3]
  PIN instruction[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END instruction[4]
  PIN instruction[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 30.640 431.580 31.240 ;
    END
  END instruction[5]
  PIN instruction[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 132.640 431.580 133.240 ;
    END
  END instruction[6]
  PIN instruction[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 438.300 110.770 442.300 ;
    END
  END instruction[7]
  PIN instruction[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 438.300 274.070 442.300 ;
    END
  END instruction[8]
  PIN instruction[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END instruction[9]
  PIN pc[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END pc[0]
  PIN pc[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 438.300 188.970 442.300 ;
    END
  END pc[10]
  PIN pc[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END pc[11]
  PIN pc[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END pc[12]
  PIN pc[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END pc[13]
  PIN pc[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END pc[14]
  PIN pc[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 234.640 431.580 235.240 ;
    END
  END pc[15]
  PIN pc[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 438.300 264.870 442.300 ;
    END
  END pc[16]
  PIN pc[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 438.300 119.970 442.300 ;
    END
  END pc[17]
  PIN pc[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END pc[18]
  PIN pc[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END pc[19]
  PIN pc[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END pc[1]
  PIN pc[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END pc[20]
  PIN pc[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END pc[21]
  PIN pc[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 438.300 292.470 442.300 ;
    END
  END pc[22]
  PIN pc[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END pc[23]
  PIN pc[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END pc[24]
  PIN pc[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END pc[25]
  PIN pc[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 438.300 101.570 442.300 ;
    END
  END pc[26]
  PIN pc[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 438.300 94.670 442.300 ;
    END
  END pc[27]
  PIN pc[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END pc[28]
  PIN pc[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END pc[29]
  PIN pc[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END pc[2]
  PIN pc[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 438.300 377.570 442.300 ;
    END
  END pc[30]
  PIN pc[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 258.440 431.580 259.040 ;
    END
  END pc[31]
  PIN pc[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END pc[3]
  PIN pc[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END pc[4]
  PIN pc[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END pc[5]
  PIN pc[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END pc[6]
  PIN pc[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 336.640 431.580 337.240 ;
    END
  END pc[7]
  PIN pc[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 81.640 431.580 82.240 ;
    END
  END pc[8]
  PIN pc[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END pc[9]
  PIN rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 438.300 25.670 442.300 ;
    END
  END rdata[0]
  PIN rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END rdata[10]
  PIN rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END rdata[11]
  PIN rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 272.040 431.580 272.640 ;
    END
  END rdata[12]
  PIN rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END rdata[13]
  PIN rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END rdata[14]
  PIN rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END rdata[15]
  PIN rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END rdata[16]
  PIN rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END rdata[17]
  PIN rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 207.440 431.580 208.040 ;
    END
  END rdata[18]
  PIN rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 438.300 179.770 442.300 ;
    END
  END rdata[19]
  PIN rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END rdata[1]
  PIN rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 438.300 205.070 442.300 ;
    END
  END rdata[20]
  PIN rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 438.300 402.870 442.300 ;
    END
  END rdata[21]
  PIN rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 425.040 431.580 425.640 ;
    END
  END rdata[22]
  PIN rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 221.040 431.580 221.640 ;
    END
  END rdata[23]
  PIN rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END rdata[24]
  PIN rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END rdata[25]
  PIN rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END rdata[26]
  PIN rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END rdata[27]
  PIN rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 193.840 431.580 194.440 ;
    END
  END rdata[28]
  PIN rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 438.300 248.770 442.300 ;
    END
  END rdata[29]
  PIN rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 295.840 431.580 296.440 ;
    END
  END rdata[2]
  PIN rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 438.300 421.270 442.300 ;
    END
  END rdata[30]
  PIN rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END rdata[31]
  PIN rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END rdata[3]
  PIN rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 146.240 431.580 146.840 ;
    END
  END rdata[4]
  PIN rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 95.240 431.580 95.840 ;
    END
  END rdata[5]
  PIN rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 438.300 129.170 442.300 ;
    END
  END rdata[6]
  PIN rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 438.300 16.470 442.300 ;
    END
  END rdata[7]
  PIN rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END rdata[8]
  PIN rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 438.300 308.570 442.300 ;
    END
  END rdata[9]
  PIN ren
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END ren
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 309.440 431.580 310.040 ;
    END
  END rst
  PIN wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END wdata[0]
  PIN wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END wdata[10]
  PIN wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 438.300 60.170 442.300 ;
    END
  END wdata[11]
  PIN wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wdata[12]
  PIN wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 438.300 395.970 442.300 ;
    END
  END wdata[13]
  PIN wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 170.040 431.580 170.640 ;
    END
  END wdata[14]
  PIN wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 438.300 239.570 442.300 ;
    END
  END wdata[15]
  PIN wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 438.300 163.670 442.300 ;
    END
  END wdata[16]
  PIN wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wdata[17]
  PIN wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END wdata[18]
  PIN wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 360.440 431.580 361.040 ;
    END
  END wdata[19]
  PIN wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 323.040 431.580 323.640 ;
    END
  END wdata[1]
  PIN wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wdata[20]
  PIN wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 438.300 326.970 442.300 ;
    END
  END wdata[21]
  PIN wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wdata[22]
  PIN wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 68.040 431.580 68.640 ;
    END
  END wdata[23]
  PIN wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 438.300 145.270 442.300 ;
    END
  END wdata[24]
  PIN wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 244.840 431.580 245.440 ;
    END
  END wdata[25]
  PIN wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 346.840 431.580 347.440 ;
    END
  END wdata[26]
  PIN wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 438.300 361.470 442.300 ;
    END
  END wdata[27]
  PIN wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 438.300 299.370 442.300 ;
    END
  END wdata[28]
  PIN wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END wdata[29]
  PIN wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wdata[2]
  PIN wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END wdata[30]
  PIN wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 438.300 223.470 442.300 ;
    END
  END wdata[31]
  PIN wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wdata[3]
  PIN wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END wdata[4]
  PIN wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 438.300 368.370 442.300 ;
    END
  END wdata[5]
  PIN wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 438.300 136.070 442.300 ;
    END
  END wdata[6]
  PIN wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 183.640 431.580 184.240 ;
    END
  END wdata[7]
  PIN wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END wdata[8]
  PIN wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 438.300 232.670 442.300 ;
    END
  END wdata[9]
  PIN wen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 54.440 431.580 55.040 ;
    END
  END wen
  PIN wstrobe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 427.580 17.040 431.580 17.640 ;
    END
  END wstrobe[0]
  PIN wstrobe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 438.300 214.270 442.300 ;
    END
  END wstrobe[1]
  PIN wstrobe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END wstrobe[2]
  PIN wstrobe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END wstrobe[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 430.000 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 430.000 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 430.000 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 425.960 334.450 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 425.960 181.270 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 425.960 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 430.000 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 430.000 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 430.000 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 425.960 411.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 425.960 257.860 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 425.960 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 8.925 425.960 429.845 ;
      LAYER met1 ;
        RECT 5.520 7.860 425.960 430.740 ;
      LAYER met2 ;
        RECT 2.390 438.020 6.710 438.300 ;
        RECT 7.550 438.020 15.910 438.300 ;
        RECT 16.750 438.020 25.110 438.300 ;
        RECT 25.950 438.020 34.310 438.300 ;
        RECT 35.150 438.020 41.210 438.300 ;
        RECT 42.050 438.020 50.410 438.300 ;
        RECT 51.250 438.020 59.610 438.300 ;
        RECT 60.450 438.020 66.510 438.300 ;
        RECT 67.350 438.020 75.710 438.300 ;
        RECT 76.550 438.020 84.910 438.300 ;
        RECT 85.750 438.020 94.110 438.300 ;
        RECT 94.950 438.020 101.010 438.300 ;
        RECT 101.850 438.020 110.210 438.300 ;
        RECT 111.050 438.020 119.410 438.300 ;
        RECT 120.250 438.020 128.610 438.300 ;
        RECT 129.450 438.020 135.510 438.300 ;
        RECT 136.350 438.020 144.710 438.300 ;
        RECT 145.550 438.020 153.910 438.300 ;
        RECT 154.750 438.020 163.110 438.300 ;
        RECT 163.950 438.020 170.010 438.300 ;
        RECT 170.850 438.020 179.210 438.300 ;
        RECT 180.050 438.020 188.410 438.300 ;
        RECT 189.250 438.020 197.610 438.300 ;
        RECT 198.450 438.020 204.510 438.300 ;
        RECT 205.350 438.020 213.710 438.300 ;
        RECT 214.550 438.020 222.910 438.300 ;
        RECT 223.750 438.020 232.110 438.300 ;
        RECT 232.950 438.020 239.010 438.300 ;
        RECT 239.850 438.020 248.210 438.300 ;
        RECT 249.050 438.020 257.410 438.300 ;
        RECT 258.250 438.020 264.310 438.300 ;
        RECT 265.150 438.020 273.510 438.300 ;
        RECT 274.350 438.020 282.710 438.300 ;
        RECT 283.550 438.020 291.910 438.300 ;
        RECT 292.750 438.020 298.810 438.300 ;
        RECT 299.650 438.020 308.010 438.300 ;
        RECT 308.850 438.020 317.210 438.300 ;
        RECT 318.050 438.020 326.410 438.300 ;
        RECT 327.250 438.020 333.310 438.300 ;
        RECT 334.150 438.020 342.510 438.300 ;
        RECT 343.350 438.020 351.710 438.300 ;
        RECT 352.550 438.020 360.910 438.300 ;
        RECT 361.750 438.020 367.810 438.300 ;
        RECT 368.650 438.020 377.010 438.300 ;
        RECT 377.850 438.020 386.210 438.300 ;
        RECT 387.050 438.020 395.410 438.300 ;
        RECT 396.250 438.020 402.310 438.300 ;
        RECT 403.150 438.020 411.510 438.300 ;
        RECT 412.350 438.020 420.710 438.300 ;
        RECT 421.550 438.020 427.610 438.300 ;
        RECT 2.390 4.280 428.100 438.020 ;
        RECT 2.950 3.555 9.010 4.280 ;
        RECT 9.850 3.555 18.210 4.280 ;
        RECT 19.050 3.555 27.410 4.280 ;
        RECT 28.250 3.555 34.310 4.280 ;
        RECT 35.150 3.555 43.510 4.280 ;
        RECT 44.350 3.555 52.710 4.280 ;
        RECT 53.550 3.555 61.910 4.280 ;
        RECT 62.750 3.555 68.810 4.280 ;
        RECT 69.650 3.555 78.010 4.280 ;
        RECT 78.850 3.555 87.210 4.280 ;
        RECT 88.050 3.555 96.410 4.280 ;
        RECT 97.250 3.555 103.310 4.280 ;
        RECT 104.150 3.555 112.510 4.280 ;
        RECT 113.350 3.555 121.710 4.280 ;
        RECT 122.550 3.555 130.910 4.280 ;
        RECT 131.750 3.555 137.810 4.280 ;
        RECT 138.650 3.555 147.010 4.280 ;
        RECT 147.850 3.555 156.210 4.280 ;
        RECT 157.050 3.555 165.410 4.280 ;
        RECT 166.250 3.555 172.310 4.280 ;
        RECT 173.150 3.555 181.510 4.280 ;
        RECT 182.350 3.555 190.710 4.280 ;
        RECT 191.550 3.555 197.610 4.280 ;
        RECT 198.450 3.555 206.810 4.280 ;
        RECT 207.650 3.555 216.010 4.280 ;
        RECT 216.850 3.555 225.210 4.280 ;
        RECT 226.050 3.555 232.110 4.280 ;
        RECT 232.950 3.555 241.310 4.280 ;
        RECT 242.150 3.555 250.510 4.280 ;
        RECT 251.350 3.555 259.710 4.280 ;
        RECT 260.550 3.555 266.610 4.280 ;
        RECT 267.450 3.555 275.810 4.280 ;
        RECT 276.650 3.555 285.010 4.280 ;
        RECT 285.850 3.555 294.210 4.280 ;
        RECT 295.050 3.555 301.110 4.280 ;
        RECT 301.950 3.555 310.310 4.280 ;
        RECT 311.150 3.555 319.510 4.280 ;
        RECT 320.350 3.555 328.710 4.280 ;
        RECT 329.550 3.555 335.610 4.280 ;
        RECT 336.450 3.555 344.810 4.280 ;
        RECT 345.650 3.555 354.010 4.280 ;
        RECT 354.850 3.555 363.210 4.280 ;
        RECT 364.050 3.555 370.110 4.280 ;
        RECT 370.950 3.555 379.310 4.280 ;
        RECT 380.150 3.555 388.510 4.280 ;
        RECT 389.350 3.555 395.410 4.280 ;
        RECT 396.250 3.555 404.610 4.280 ;
        RECT 405.450 3.555 413.810 4.280 ;
        RECT 414.650 3.555 423.010 4.280 ;
        RECT 423.850 3.555 428.100 4.280 ;
      LAYER met3 ;
        RECT 4.400 434.840 427.580 435.705 ;
        RECT 2.365 426.040 427.580 434.840 ;
        RECT 2.365 424.640 427.180 426.040 ;
        RECT 2.365 422.640 427.580 424.640 ;
        RECT 4.400 421.240 427.580 422.640 ;
        RECT 2.365 412.440 427.580 421.240 ;
        RECT 2.365 411.040 427.180 412.440 ;
        RECT 2.365 409.040 427.580 411.040 ;
        RECT 4.400 407.640 427.580 409.040 ;
        RECT 2.365 398.840 427.580 407.640 ;
        RECT 2.365 397.440 427.180 398.840 ;
        RECT 2.365 395.440 427.580 397.440 ;
        RECT 4.400 394.040 427.580 395.440 ;
        RECT 2.365 388.640 427.580 394.040 ;
        RECT 2.365 387.240 427.180 388.640 ;
        RECT 2.365 385.240 427.580 387.240 ;
        RECT 4.400 383.840 427.580 385.240 ;
        RECT 2.365 375.040 427.580 383.840 ;
        RECT 2.365 373.640 427.180 375.040 ;
        RECT 2.365 371.640 427.580 373.640 ;
        RECT 4.400 370.240 427.580 371.640 ;
        RECT 2.365 361.440 427.580 370.240 ;
        RECT 2.365 360.040 427.180 361.440 ;
        RECT 2.365 358.040 427.580 360.040 ;
        RECT 4.400 356.640 427.580 358.040 ;
        RECT 2.365 347.840 427.580 356.640 ;
        RECT 2.365 346.440 427.180 347.840 ;
        RECT 2.365 344.440 427.580 346.440 ;
        RECT 4.400 343.040 427.580 344.440 ;
        RECT 2.365 337.640 427.580 343.040 ;
        RECT 2.365 336.240 427.180 337.640 ;
        RECT 2.365 334.240 427.580 336.240 ;
        RECT 4.400 332.840 427.580 334.240 ;
        RECT 2.365 324.040 427.580 332.840 ;
        RECT 2.365 322.640 427.180 324.040 ;
        RECT 2.365 320.640 427.580 322.640 ;
        RECT 4.400 319.240 427.580 320.640 ;
        RECT 2.365 310.440 427.580 319.240 ;
        RECT 2.365 309.040 427.180 310.440 ;
        RECT 2.365 307.040 427.580 309.040 ;
        RECT 4.400 305.640 427.580 307.040 ;
        RECT 2.365 296.840 427.580 305.640 ;
        RECT 2.365 295.440 427.180 296.840 ;
        RECT 2.365 293.440 427.580 295.440 ;
        RECT 4.400 292.040 427.580 293.440 ;
        RECT 2.365 286.640 427.580 292.040 ;
        RECT 2.365 285.240 427.180 286.640 ;
        RECT 2.365 283.240 427.580 285.240 ;
        RECT 4.400 281.840 427.580 283.240 ;
        RECT 2.365 273.040 427.580 281.840 ;
        RECT 2.365 271.640 427.180 273.040 ;
        RECT 2.365 269.640 427.580 271.640 ;
        RECT 4.400 268.240 427.580 269.640 ;
        RECT 2.365 259.440 427.580 268.240 ;
        RECT 2.365 258.040 427.180 259.440 ;
        RECT 2.365 256.040 427.580 258.040 ;
        RECT 4.400 254.640 427.580 256.040 ;
        RECT 2.365 245.840 427.580 254.640 ;
        RECT 4.400 244.440 427.180 245.840 ;
        RECT 2.365 235.640 427.580 244.440 ;
        RECT 2.365 234.240 427.180 235.640 ;
        RECT 2.365 232.240 427.580 234.240 ;
        RECT 4.400 230.840 427.580 232.240 ;
        RECT 2.365 222.040 427.580 230.840 ;
        RECT 2.365 220.640 427.180 222.040 ;
        RECT 2.365 218.640 427.580 220.640 ;
        RECT 4.400 217.240 427.580 218.640 ;
        RECT 2.365 208.440 427.580 217.240 ;
        RECT 2.365 207.040 427.180 208.440 ;
        RECT 2.365 205.040 427.580 207.040 ;
        RECT 4.400 203.640 427.580 205.040 ;
        RECT 2.365 194.840 427.580 203.640 ;
        RECT 4.400 193.440 427.180 194.840 ;
        RECT 2.365 184.640 427.580 193.440 ;
        RECT 2.365 183.240 427.180 184.640 ;
        RECT 2.365 181.240 427.580 183.240 ;
        RECT 4.400 179.840 427.580 181.240 ;
        RECT 2.365 171.040 427.580 179.840 ;
        RECT 2.365 169.640 427.180 171.040 ;
        RECT 2.365 167.640 427.580 169.640 ;
        RECT 4.400 166.240 427.580 167.640 ;
        RECT 2.365 157.440 427.580 166.240 ;
        RECT 2.365 156.040 427.180 157.440 ;
        RECT 2.365 154.040 427.580 156.040 ;
        RECT 4.400 152.640 427.580 154.040 ;
        RECT 2.365 147.240 427.580 152.640 ;
        RECT 2.365 145.840 427.180 147.240 ;
        RECT 2.365 143.840 427.580 145.840 ;
        RECT 4.400 142.440 427.580 143.840 ;
        RECT 2.365 133.640 427.580 142.440 ;
        RECT 2.365 132.240 427.180 133.640 ;
        RECT 2.365 130.240 427.580 132.240 ;
        RECT 4.400 128.840 427.580 130.240 ;
        RECT 2.365 120.040 427.580 128.840 ;
        RECT 2.365 118.640 427.180 120.040 ;
        RECT 2.365 116.640 427.580 118.640 ;
        RECT 4.400 115.240 427.580 116.640 ;
        RECT 2.365 106.440 427.580 115.240 ;
        RECT 2.365 105.040 427.180 106.440 ;
        RECT 2.365 103.040 427.580 105.040 ;
        RECT 4.400 101.640 427.580 103.040 ;
        RECT 2.365 96.240 427.580 101.640 ;
        RECT 2.365 94.840 427.180 96.240 ;
        RECT 2.365 92.840 427.580 94.840 ;
        RECT 4.400 91.440 427.580 92.840 ;
        RECT 2.365 82.640 427.580 91.440 ;
        RECT 2.365 81.240 427.180 82.640 ;
        RECT 2.365 79.240 427.580 81.240 ;
        RECT 4.400 77.840 427.580 79.240 ;
        RECT 2.365 69.040 427.580 77.840 ;
        RECT 2.365 67.640 427.180 69.040 ;
        RECT 2.365 65.640 427.580 67.640 ;
        RECT 4.400 64.240 427.580 65.640 ;
        RECT 2.365 55.440 427.580 64.240 ;
        RECT 2.365 54.040 427.180 55.440 ;
        RECT 2.365 52.040 427.580 54.040 ;
        RECT 4.400 50.640 427.580 52.040 ;
        RECT 2.365 45.240 427.580 50.640 ;
        RECT 2.365 43.840 427.180 45.240 ;
        RECT 2.365 41.840 427.580 43.840 ;
        RECT 4.400 40.440 427.580 41.840 ;
        RECT 2.365 31.640 427.580 40.440 ;
        RECT 2.365 30.240 427.180 31.640 ;
        RECT 2.365 28.240 427.580 30.240 ;
        RECT 4.400 26.840 427.580 28.240 ;
        RECT 2.365 18.040 427.580 26.840 ;
        RECT 2.365 16.640 427.180 18.040 ;
        RECT 2.365 14.640 427.580 16.640 ;
        RECT 4.400 13.240 427.580 14.640 ;
        RECT 2.365 4.440 427.580 13.240 ;
        RECT 2.365 3.575 427.180 4.440 ;
      LAYER met4 ;
        RECT 9.070 13.095 20.640 428.225 ;
        RECT 23.040 13.095 97.440 428.225 ;
        RECT 99.840 13.095 174.240 428.225 ;
        RECT 176.640 13.095 251.040 428.225 ;
        RECT 253.440 13.095 327.840 428.225 ;
        RECT 330.240 13.095 404.640 428.225 ;
        RECT 407.040 13.095 412.785 428.225 ;
      LAYER met5 ;
        RECT 8.860 182.870 393.180 240.500 ;
        RECT 8.860 106.280 393.180 178.070 ;
        RECT 8.860 29.690 393.180 101.480 ;
        RECT 8.860 17.900 393.180 24.890 ;
  END
END core
END LIBRARY

