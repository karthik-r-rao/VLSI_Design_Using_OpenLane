
.SUBCKT sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z net35 sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net39 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net39 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net35 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB net35 Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net39 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net35 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_8 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_2 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_1 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_4 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkinvkapwr_16 A KAPWR VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A KAPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net87 net153 net117 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net117 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net110 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net98 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net98 M1 net110 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net153 clkneg net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net87 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net93 net87 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net153 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net87 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net87 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net153 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net87 net153 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net87 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net153 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B majb VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs1 sumb majb nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs20 VGND A nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs21 VGND B nint1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 majb A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 majb B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1 VPWR majb sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs20 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs21 sndPA B sumb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net82 s0 net108 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net101 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net93 M1 net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net82 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net81 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net165 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net82 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net165 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net82 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net144 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net82 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=1 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
MI36 net120 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net103 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net71 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net120 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net88 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net80 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net80 S1 net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net71 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net103 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net128 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net128 VGND VNB nfet_01v8 m=5 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net179 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net179 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net156 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net143 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net143 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net128 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net128 VPWR VPB pfet_01v8_hvt m=5 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net125 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
rI12 VGND LO short
rI11 HI VPWR short
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net138 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net78 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net78 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net54 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net54 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 net163 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net163 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net195 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net195 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net130 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net130 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net107 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI34 S0 clkpos net219 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net239 S1 net187 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net230 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net199 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net230 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net219 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net239 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net199 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net195 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net187 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net195 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net159 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net159 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net138 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net138 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net199 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net199 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net98 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net98 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI27 net243 S1 net215 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net230 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net227 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net199 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net215 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net206 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net199 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net227 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net230 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net243 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net83 net121 net109 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net109 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net102 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net94 M1 net102 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net121 clkneg net82 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net83 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net82 net83 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos net121 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net166 net83 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net83 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 net121 clkpos net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net83 net121 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net145 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net145 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net145 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net83 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg net121 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_2 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_1 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__maj3_4 A B C VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net55 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net55 net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 X net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net55 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net55 net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 X net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net104 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net104 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net189 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net169 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net189 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net169 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
MI645 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net165 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net165 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net96 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkpos net96 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net84 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net84 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net212 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net209 S1 net157 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net200 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net196 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net212 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net209 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net196 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net165 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net157 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net165 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_8 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_4 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_16 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_2 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_clkbufkapwr_1 A KAPWR VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab KAPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
MI1 VGND VPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 VPWR VGND VPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd2_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 A LOWLVPWR VGND VPB VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 A LOWLVPWR VGND VPB VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A LOWLVPWR LOWLVPWR pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_4 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.05 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.05 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_8 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=2.89 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=2.89 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_12 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=4.73 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=4.73 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_6 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=1.97 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=1.97 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_decapkapwr_3 KAPWR VGND VNB VPB VPWR
MI1 VGND KAPWR VGND VNB nfet_01v8 m=1 w=0.55 l=0.59 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 KAPWR VGND KAPWR VPB pfet_01v8_hvt m=1 w=0.87 l=0.59 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
MMNA00 xb A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 xb A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X xb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 xb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X xb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net92 S0 net134 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net134 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net127 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net115 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net115 M1 net127 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net103 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net92 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net103 net92 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI672 net171 net92 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 Q_N net171 VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net215 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net92 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net215 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net92 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net194 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net92 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI673 net171 net92 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI671 Q_N net171 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
MMNA00 Y A0 smdNA0 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 sndNA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S sndPS VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb sndPSb VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_1 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_4 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor3_2 A B C VGND VNB VPB VPWR X
MMIP3 X net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 Cb net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 mid2 C net117 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 C net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 Cb net117 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1p_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA A net36 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 VPWR net36 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net36 SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net121 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net121 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net125 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net61 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net125 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net61 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net57 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net57 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net125 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net125 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net108 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net116 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net116 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net108 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net96 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 pndA A4 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 sndA3 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 sndA3 A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
MI662 net88 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net88 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net76 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net76 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 net63 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 net116 GATE net63 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net76 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net116 clkneg M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net116 clkpos M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net123 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net123 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 net116 SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net76 m1 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net116 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net76 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 A LOWLVPWR VGND VNB VPB VPWR X
MI2 net72 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 cross1 net72 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Ab A LOWLVPWR LOWLVPWR pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 X net60 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 net60 cross1 VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 cross1 Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net72 A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 X net60 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 net60 cross1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0n_1 A SLEEP_B VGND VNB VPB VPWR X
MI14 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net36 A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 sndA SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 net36 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 Y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_2 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_1 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_4 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_0 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA net25 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net25 TE_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net25 TE_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvn_8 A TE_B VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TE TE_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TE_B sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TE TE_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s6s_1 A VGND VNB VPB VPWR X
MMIN1 Ab net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net56 net48 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net52 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net48 net44 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net44 net52 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net56 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net56 net48 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net48 net44 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net44 net52 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net52 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s18_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__probe_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net29 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net29 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net29 X short
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
MMIN0 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
MMNA00 sndNS0ba0 S0b xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 sndNS0ba0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 xlowb VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 sndNS0a1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 sndNS0ba2 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 xhib VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 sndNS0a3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b xlowb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 xhib VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 S1b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 S0b VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 sndPA0a0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b sndPA1a1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 sndPA2a2 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b sndPA3a3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 xlowb VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMPs2o xb S1b xhib VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 S1b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 S0b VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.028 perim=0.76
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=24 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=8 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
MMIN0 Y A VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 A VGND VPB VPWRIN VPWR X
M1000 X a_1028_32# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.1725e+11p pd=2.13e+06u as=4.7795e+11p ps=4.37e+06u
M1001 VPWR a_620_911# a_714_58# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
M1002 a_1028_32# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1003 X a_1028_32# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.8525e+11p pd=1.87e+06u as=1.4178e+12p ps=1.319e+07u
M1004 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=0p ps=0u
M1005 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1006 a_714_58# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1007 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1008 a_1028_32# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1009 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1010 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1012 VGND A a_714_58# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1014 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_714_58# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=1.1152e+12p pd=9.97e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u
+ ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1003 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.81105e+12p ps=1.7e+07u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1005 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1006 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=4.225e+11p pd=3.9e+06u as=0p ps=0u
M1007 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1008 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1009 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1010 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1011 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1012 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1013 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1014 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1015 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1016 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1017 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1018 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1019 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1020 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 A VGND VPB VPWRIN VPWR X
M1000 VPWR a_620_911# a_714_47# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=8.352e+11p pd=7.41e+06u as=2.1725e+11p ps=2.13e+06u
M1001 a_1032_911# a_620_911# VPWR VPB pfet_01v8_hvt w=790000u
+ l=150000u ad=2.133e+11p pd=2.12e+06u as=0p ps=0u
M1002 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=3.64e+11p pd=3.72e+06u as=1.62905e+12p ps=1.514e+07u
M1003 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=3.64e+11p
+ pd=3.72e+06u as=0p ps=0u
M1004 a_714_47# A VGND VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1005 X a_1032_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=2.405e+11p pd=2.04e+06u as=0p ps=0u
M1006 VPWR a_1032_911# X VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=3.7e+11p ps=2.74e+06u
M1007 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1008 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1009 a_1032_911# a_620_911# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1010 VGND A a_714_47# VGND nfet_01v8 w=650000u l=150000u ad=0p pd=0u
+ as=0p ps=0u
M1011 a_505_297# A VPWRIN VPWRIN pfet_01v8_hvt w=1e+06u l=150000u
+ ad=2.75e+11p pd=2.55e+06u as=2.75e+11p ps=2.55e+06u
M1012 a_505_297# A VGND VGND nfet_01v8 w=420000u l=150000u
+ ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 X a_1032_911# VPWR VPB pfet_01v8_hvt w=1e+06u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1014 VGND a_1032_911# X VGND nfet_01v8 w=650000u l=150000u ad=0p
+ pd=0u as=0p ps=0u
M1015 VGND a_505_297# a_620_911# VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1016 a_620_911# a_505_297# VGND VGND nfet_01v8 w=650000u l=150000u
+ ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_714_47# a_620_911# VPB pfet_01v8_hvt w=790000u l=150000u
+ ad=0p pd=0u as=2.1725e+11p ps=2.13e+06u
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMIP3 SUM net144 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bbb Bb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CINb1 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CINbb2 CINb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CINb2 CIN VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CINbb2 mid2 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CINb2 mid1 net144 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bbb mid2 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CINb1 mid1 COUT VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net144 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CINb1 mid2 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CINb1 CIN VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CINbb2 CINb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CINb2 CIN VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CINbb2 mid1 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CINb2 mid2 net144 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bbb mid1 COUT VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bbb Bb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_2 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__probec_p_8 A VGND VNB VPB VPWR X
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net33 Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net33 Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
rI112 net33 X short
rI120 VGND met5vgnd short
rI119 VPWR met5vpwr short
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
MMIN1 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_4 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_2 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA Ab X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_16 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrc_8 A SLEEP VGND VNB VPB VPWR X
MMP0 VPWR Ab sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA SLEEP X VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 X SLEEP VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_bleeder_1 SHORT VGND VNB VPB VPWR
MI2 net29 SHORT net25 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net25 SHORT net24 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 VPWR SHORT net29 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 net24 SHORT net16 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net16 SHORT VGND VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_2 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net128 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net111 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net96 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net88 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net88 S1 net96 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net111 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net140 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net140 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net191 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net191 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net168 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net168 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net155 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net140 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net140 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
MI36 net129 M0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M1 M0 net112 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net80 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 S0 clkpos net129 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net97 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 S0 clkneg net89 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 net89 S1 net97 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 S1 S0 VGND VNB nfet_01v8 m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkpos net80 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net112 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net141 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net141 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 Q_N S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 S0 clkneg net192 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net192 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net156 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 S0 clkpos net156 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 S0 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net141 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net141 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
MMNnand0 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA B inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 y inand nmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 y inand VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlygate4sd2_1 A VGND VNB VPB VPWR X
MMIN1 Ab net34 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net34 net30 VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net30 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab net34 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net34 net30 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net30 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=12 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=12 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=1 w=0.52 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=1 w=0.79 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X Ab VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj31 sndNCINn3 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND A sndNCINn3 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR A sndPCINp3 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 sndPCINp3 CIN majb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj31 sndPCINp3 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
MMNs1s nint1 majb sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 COUT majb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM sumb VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj10 majb B sndNAp1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj11 sndNAp1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj30 majb CIN nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj21 nmajmid A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNmaj20 VGND B nmajmid VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s0 VGND A sndNAn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s1 sndNAn4 B sndNBn4 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs2s2 sndNBn4 CIN sumb VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s0 nint1 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s1 nint1 B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNs3s2 nint1 CIN VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT majb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM sumb VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj10 VPWR A sndPAp1 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj11 sndPAp1 B majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj20 VPWR B pmajmid VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj30 pmajmid CIN majb VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPmaj21 pmajmid A VPWR VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s0 VPWR A sndPAp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s1 sndPAp4 B sndPBp4 VPB pfet_01v8_hvt m=1 w=0.63 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs2s2 sndPBp4 CIN sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s0 pint1 A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s1 pint1 B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs3s2 pint1 CIN VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPs1s pint1 majb sumb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbn_1 D GATE_N VGND VNB VPB VPWR Q Q_N
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net112 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net56 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net112 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net56 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net52 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net52 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net112 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net112 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net107 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net107 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net87 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net87 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_0 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.7 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_8 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
MMIN1 Ab A VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Y Abb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 Y Abb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 A SLEEP KAPWR VGND VNB VPB VPWR X
MMP0 VPWR SLEEP sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA net58 net66 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 net58 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 Ab net66 KAPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 X Ab KAPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net66 SLEEP VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 net66 net58 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 net58 A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Ab net66 VGND VNB nfet_01v8 m=4 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 X Ab VGND VNB nfet_01v8 m=16 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 pndB B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_0 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
MMPA0 net40 A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 net40 A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 net40 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net123 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net123 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net235 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net235 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net203 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net203 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
MI14 net155 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net155 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net144 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net127 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net127 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net144 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net116 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net107 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net104 D net116 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net104 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net104 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 Q_N q1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net240 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net240 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net224 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net224 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net104 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net104 D net180 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net200 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net200 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net192 q1 net104 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net192 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net180 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net176 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net176 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 Q_N q1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 Q_N net114 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net58 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 net114 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkneg GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net58 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net54 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkneg GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 Q_N net114 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 net114 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net109 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net109 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net89 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net89 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
MMIP3 SUM net146 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 Bb2 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab Bb1 mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb Bb1 mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 CIb1 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 CIbb2 CIb2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 CIb2 CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb1 B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb2 mid2 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb2 mid1 net146 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb2 mid2 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb1 mid1 COUT_N VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net146 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb1 mid2 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb Bb1 mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab Bb1 mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 CIb1 CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 CIbb2 CIb2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 CIb2 CI VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb1 B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb2 mid1 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb2 mid2 net146 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 Bb2 mid1 COUT_N VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Bb2 B VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net190 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net190 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net99 s0 net125 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net125 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net118 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net110 M1 net118 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net98 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net99 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net98 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI53 net142 net99 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI50 Q_N net142 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net181 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net99 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net181 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net99 s0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net169 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net169 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net169 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net99 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI52 net142 net99 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI51 Q_N net142 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_16 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=6 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=16 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=16 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=6 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__bufbuf_8 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 Abb Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 Abbb Abb VGND VNB nfet_01v8 m=3 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X Abbb VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X Abbb VPWR VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Abbb Abb VPWR VPB pfet_01v8_hvt m=3 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputisolatch_1 D SLEEP_B VGND VNB VPB VPWR Q
MI677 Q s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 sleepneg sleeppos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI674 net39 s0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 s0 sleepneg net49 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net49 D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 sleeppos net38 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net38 net39 VGND VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 sleeppos SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 sleeppos SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 sleepneg sleeppos VPWR VPB pfet_01v8_hvt m=1 w=0.55 l=0.15
+ mult=1 sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063
+ perim=1.14
MI662 net86 net39 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 sleepneg net86 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net39 s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q s0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 s0 sleeppos net69 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net69 D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_4 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=4 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=8 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=8 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=8 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_1 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
MMN0 Z A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA TE VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 TEB TE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR TEB sndTEB VPB pfet_01v8_hvt m=2 w=0.94 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndTEB A Z VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 TEB TE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 VPWR D1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 pndC C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 pndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
MI657 M0 clkpos net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net96 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 net88 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net72 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net72 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 Q_N net88 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net128 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net147 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net88 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net147 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net128 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 Q_N net88 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
MI14 net115 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net115 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net59 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net79 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net83 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net83 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net79 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net76 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net76 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net59 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net175 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net175 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net172 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net160 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net148 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net148 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net172 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net128 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net128 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
MMNnor0 inor A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND A sndNA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNA B X VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 X inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA B inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 X inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
MMIN1 Ab X VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 net59 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X net47 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 net51 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net47 net43 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net43 net51 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab X VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 net59 Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 X net47 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 net47 net43 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net43 net51 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 net51 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
MI662 net75 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M0 clkpos net75 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net63 CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net63 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 net54 GATE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 GCLK net63 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 M0 clkneg net110 VNB nfet_01v8 m=1 w=0.39 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 M0 clkpos net91 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net99 CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net63 m1 net99 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 net91 GATE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 GCLK net63 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnand0 VGND A1_N sndNA1N VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnand1 sndNA1N A2_N inand VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 nmid B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 nmid B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inand nmid VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand0 inand A1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnand1 inand A2_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 VPWR B1 sndPB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 sndPB1 B2 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inand VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
MMIN2 COUT net195 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 SUM net123 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 CIb mid2 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Bb mid1 net195 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 CIbb mid2 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 CIb mid1 net123 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 CIbb CIb VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 CIb CI VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Ab2 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 Abb2 Ab2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI14 Ab1 A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 Abb2 B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Ab1 Bb mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Abb2 Bb mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Ab1 B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 COUT net195 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 SUM net123 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 CIb mid1 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 Bb mid2 net195 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI1 CIbb mid1 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 CIb mid2 net123 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 CIbb CIb VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 CIb CI VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 Ab2 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 Abb2 Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 Ab1 A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Abb2 Bb mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 Ab1 B mid1 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 Abb2 B mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 Ab1 Bb mid2 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
MI14 net124 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net124 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 net68 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net109 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net92 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net92 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net109 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net85 DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 db S1 net85 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 db D net68 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 Q_N S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net193 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net193 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net148 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net168 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net168 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 S1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net161 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net161 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 db D net148 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 db S1 net141 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI12 net141 deneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI22 Q_N S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 VPWR C1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 pndB B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 pndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net90 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net90 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
MI642 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net84 S0 net114 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net114 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net95 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net95 M1 net107 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net83 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 Q net84 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net83 net84 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net187 net84 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net84 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net187 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net84 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net166 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net166 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net166 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 Q net84 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.54 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_0 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 sndB1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 y B2 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso0p_1 A SLEEP VGND VNB VPB VPWR X
MI8 net36 A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net36 sleepb VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 X net36 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 sleepb SLEEP VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net36 sleepb sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI21 X net36 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 sleepb SLEEP VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 sndA A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__tap_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 D D_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 Y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 D D_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 Y B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 Y C VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPB1N B1 B1_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINB1N B1 B1_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net55 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net55 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net51 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net94 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net102 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net102 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net94 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net82 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net82 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net54 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 m1 RESET_B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net54 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net50 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net50 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net93 RESET_B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net101 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net101 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 net93 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net81 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net81 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2111oi_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 pndC C1 pndB VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPD0 Y D1 pndC VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMND0 Y D1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_4 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_2 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__xnor3_1 A B C VGND VNB VPB VPWR X
MMIN3 X net57 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI29 Ab Bb mid2 VNB nfet_01v8 m=1 w=0.6 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 Abb Bb mid1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 Bb B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 mid1 Cb net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 Ab A VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 Cb C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI2 mid2 C net57 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 Abb Ab VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI24 Ab B mid1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI28 Abb B mid2 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X net57 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 mid1 C net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI27 mid2 B Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 Abb Ab VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 mid1 B Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI26 mid2 Bb Abb VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 mid2 Cb net57 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 Cb C VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 Bb B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 mid1 Bb Ab VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
MI657 M0 clkpos net79 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net79 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net59 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net59 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net107 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net122 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net122 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net107 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__tapvgnd_1 VGND VPB VPWR
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_2 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=2 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkdlybuf4s15_1 A VGND VNB VPB VPWR X
MMIN1 Ab A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 A2 Ab VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Ab2 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 X Ab2 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 A2 Ab VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 Ab2 A2 VPWR VPB pfet_01v8_hvt m=1 w=0.82 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 X Ab2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 Y VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 pndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
MMP0 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B sndPB VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C sndPC VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 sndPC D y VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP4 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 y D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN4 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 net36 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net36 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
MMIP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.25 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 Y A net31 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net35 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net31 A VGND VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI5 Y A net35 VNB nfet_01v8 m=1 w=0.55 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net114 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net114 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net94 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net103 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net103 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net94 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net222 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net222 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net211 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net211 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net167 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net179 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net179 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net167 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net158 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net158 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
MI14 net146 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg net146 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net135 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net118 q1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net118 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net135 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net107 deneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net98 sceneg db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD net98 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net95 D net107 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net95 SCE db VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net87 q1 net95 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE net87 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net227 q1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net227 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net206 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos net206 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net95 sceneg db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net95 D net190 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net187 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos net187 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net174 q1 net95 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg net174 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net190 DE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net163 SCE db VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD net163 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 Y C2 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 net62 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net62 C2 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 pndB B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 pndB B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPC0 Y C1 pndB VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNC0 Y C1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net53 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net53 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net44 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net96 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net96 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net76 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net76 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
MI635 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI17 M0 clkneg net51 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 Q m1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 clkpos GATE_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 net51 db VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 net47 m1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 M0 clkpos net47 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 m1 M0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 db D VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 clkpos GATE_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 Q m1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M0 clkneg net94 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net94 m1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 m1 M0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI19 M0 clkpos net74 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI20 net74 db VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 Y C VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP3 Y D VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 B B_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B sndB VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C sndC VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN3 sndC D VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 B B_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
MMP0 Y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 Y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 Y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X
MMP0 y A VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 X y VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A sndA VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 sndA B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 X y VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
MMNnor0 inor A1_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNnor1 inor A2_N VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi10 VGND B1 sndNB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi11 sndNB1 B2 Y VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNaoi20 Y inor VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor0 VPWR A1_N sndPA1N VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPnor1 sndPA1N A2_N inor VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi10 pmid B1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi11 pmid B2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPaoi20 Y inor pmid VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
MMPA0 pndA A1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 pndA A2 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 pndA A3 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 Y B1 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB1 Y B2 pndA VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 Y A1 sndA1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 sndA1 A2 sndA2 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 sndA2 A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 Y B1 sndB1 VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB1 sndB1 B2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__macro_sparecell VGND VNB VPB VPWR LO
XI1 net59 LO VGND VNB VPB VPWR / sky130_fd_sc_hd__conb_1
XI6 nor2right invright VGND VNB VPB VPWR / sky130_fd_sc_hd__inv_2
XI7 nor2left invleft VGND VNB VPB VPWR / sky130_fd_sc_hd__inv_2
XI4 nd2right nd2right nor2right VGND VNB VPB VPWR /
+ sky130_fd_sc_hd__nor2_2
XI5 nd2left nd2left nor2left VGND VNB VPB VPWR /
+ sky130_fd_sc_hd__nor2_2
XI2 LO LO nd2right VGND VNB VPB VPWR / sky130_fd_sc_hd__nand2_2
XI3 LO LO nd2left VGND VNB VPB VPWR / sky130_fd_sc_hd__nand2_2
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=4 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=4 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
MMPA0 VPWR A1 sndA1 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 sndA2 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA2 sndA2 A3 sndA3 VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA3 sndA3 A4 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 y VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA2 pndA A3 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA3 pndA A4 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 pndA VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMINX X y VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net160 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net160 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net128 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net128 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
MI98 net105 D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 net105 SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI46 clkneg clkpos VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net176 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net213 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net176 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net153 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkpos CLK_N VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net153 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net145 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net145 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net117 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net213 net117 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net105 clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net125 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net125 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net117 RESET net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net117 S0 net116 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net116 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 net105 D p0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 net105 sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net265 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net213 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net117 S0 net268 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net265 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net216 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net257 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net257 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net117 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net268 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net241 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net105 clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net241 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkneg clkpos VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkpos CLK_N VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net216 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net213 net117 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net117 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
MI46 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 db D VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 RESET RESET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI676 M1 M0 net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI675 net141 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net162 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI677 M1 RESET net141 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M0 clkpos net118 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI44 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 net118 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 S0 clkneg net110 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net110 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 Q_N net82 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net162 net82 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI668 S0 clkpos net93 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI667 net93 M1 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI630 net82 RESET net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI3 net82 S0 net81 VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 net81 SET_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI679 M1 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI669 S0 clkneg net218 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net162 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net82 S0 net221 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI670 net218 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI678 net165 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 S0 clkpos net210 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI10 net82 SET_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI11 net221 RESET VPWR VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 net194 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db D VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 M0 clkneg net194 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 RESET RESET_B VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI45 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI680 M1 M0 net165 VPB pfet_01v8_hvt m=1 w=0.84 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net162 net82 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net82 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__lpflow_inputiso1n_1 A SLEEP_B VGND VNB VPB VPWR X
MI23 VPWR A sndPA VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI8 VPWR net44 X VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 net56 SLEEP_B VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI7 sndPA net56 net44 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 net56 SLEEP_B VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI25 net44 A VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 X net44 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI9 net44 net56 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=2 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net196 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net189 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=2 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net196 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net189 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS




.SUBCKT sky130_fd_sc_hd__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
MI98 db D n0 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI657 M0 clkpos net129 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net129 M1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net120 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg net120 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S1 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg M0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI639 sceb SCE VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 M1 clkpos S0 VNB nfet_01v8 m=1 w=0.36 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N net153 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net153 S1 VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 S1 S0 VGND VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VGND VNB nfet_01v8 m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VGND VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 S1 S0 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos net177 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 M1 M0 VPWR VPB pfet_01v8_hvt m=1 w=0.75 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net160 M1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S1 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N net153 VPWR VPB pfet_01v8_hvt m=1 w=1.0 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net177 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos M0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 M1 clkneg S0 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI640 sceb SCE VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg net160 VPB pfet_01v8_hvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 net153 S1 VPWR VPB pfet_01v8_hvt m=1 w=0.64 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS






















































































































.subckt core clk data_address[0] data_address[10] data_address[11] data_address[12]
+ data_address[13] data_address[14] data_address[15] data_address[16] data_address[17]
+ data_address[18] data_address[19] data_address[1] data_address[20] data_address[21]
+ data_address[22] data_address[23] data_address[24] data_address[25] data_address[26]
+ data_address[27] data_address[28] data_address[29] data_address[2] data_address[30]
+ data_address[31] data_address[3] data_address[4] data_address[5] data_address[6]
+ data_address[7] data_address[8] data_address[9] instruction[0] instruction[10] instruction[11]
+ instruction[12] instruction[13] instruction[14] instruction[15] instruction[16]
+ instruction[17] instruction[18] instruction[19] instruction[1] instruction[20] instruction[21]
+ instruction[22] instruction[23] instruction[24] instruction[25] instruction[26]
+ instruction[27] instruction[28] instruction[29] instruction[2] instruction[30] instruction[31]
+ instruction[3] instruction[4] instruction[5] instruction[6] instruction[7] instruction[8]
+ instruction[9] pc[0] pc[10] pc[11] pc[12] pc[13] pc[14] pc[15] pc[16] pc[17] pc[18]
+ pc[19] pc[1] pc[20] pc[21] pc[22] pc[23] pc[24] pc[25] pc[26] pc[27] pc[28] pc[29]
+ pc[2] pc[30] pc[31] pc[3] pc[4] pc[5] pc[6] pc[7] pc[8] pc[9] rdata[0] rdata[10]
+ rdata[11] rdata[12] rdata[13] rdata[14] rdata[15] rdata[16] rdata[17] rdata[18]
+ rdata[19] rdata[1] rdata[20] rdata[21] rdata[22] rdata[23] rdata[24] rdata[25] rdata[26]
+ rdata[27] rdata[28] rdata[29] rdata[2] rdata[30] rdata[31] rdata[3] rdata[4] rdata[5]
+ rdata[6] rdata[7] rdata[8] rdata[9] ren rst wdata[0] wdata[10] wdata[11] wdata[12]
+ wdata[13] wdata[14] wdata[15] wdata[16] wdata[17] wdata[18] wdata[19] wdata[1] wdata[20]
+ wdata[21] wdata[22] wdata[23] wdata[24] wdata[25] wdata[26] wdata[27] wdata[28]
+ wdata[29] wdata[2] wdata[30] wdata[31] wdata[3] wdata[4] wdata[5] wdata[6] wdata[7]
+ wdata[8] wdata[9] wen wstrobe[0] wstrobe[1] wstrobe[2] wstrobe[3] VPWR VGND
X_09671_ _10808_/A VGND VGND VPWR VPWR _10415_/A sky130_fd_sc_hd__buf_1
XFILLER_27_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08622_ _08622_/A VGND VGND VPWR VPWR _08622_/X sky130_fd_sc_hd__clkbuf_1
X_08553_ _08563_/A VGND VGND VPWR VPWR _08566_/A sky130_fd_sc_hd__inv_2
XFILLER_51_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07504_ _07506_/A _12563_/A VGND VGND VPWR VPWR _15520_/D sky130_fd_sc_hd__nor2_1
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08484_ _10781_/A VGND VGND VPWR VPWR _09250_/A sky130_fd_sc_hd__buf_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07435_ _07443_/A VGND VGND VPWR VPWR _07438_/A sky130_fd_sc_hd__clkbuf_1
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07366_ _07366_/A VGND VGND VPWR VPWR _12573_/A sky130_fd_sc_hd__buf_1
X_09105_ _09105_/A VGND VGND VPWR VPWR _09105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07297_ _07297_/A VGND VGND VPWR VPWR _07363_/A sky130_fd_sc_hd__buf_1
XFILLER_148_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09036_ _09038_/A VGND VGND VPWR VPWR _09036_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09938_ _10308_/A VGND VGND VPWR VPWR _09938_/X sky130_fd_sc_hd__buf_1
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09869_ _09878_/A VGND VGND VPWR VPWR _09869_/X sky130_fd_sc_hd__buf_1
XFILLER_93_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11900_ _11900_/A VGND VGND VPWR VPWR _11905_/A sky130_fd_sc_hd__clkbuf_2
X_12880_ _13343_/X _12741_/X _12810_/A _12878_/X _12879_/Y VGND VGND VPWR VPWR _12880_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_202 _13574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_213 _13476_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11831_ _11837_/A VGND VGND VPWR VPWR _11831_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_224 _11559_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_235 _09847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_246 _11895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_257 _12651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14550_ _11486_/X _14550_/D VGND VGND VPWR VPWR _14550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11762_ _11762_/A VGND VGND VPWR VPWR _11762_/X sky130_fd_sc_hd__clkbuf_1
X_13501_ _13500_/X rdata[7] _13516_/S VGND VGND VPWR VPWR _13501_/X sky130_fd_sc_hd__mux2_2
X_10713_ _11471_/A VGND VGND VPWR VPWR _10713_/X sky130_fd_sc_hd__buf_1
X_14481_ _11749_/X _14481_/D VGND VGND VPWR VPWR _14481_/Q sky130_fd_sc_hd__dfxtp_1
X_11693_ _11725_/A VGND VGND VPWR VPWR _11716_/A sky130_fd_sc_hd__buf_2
X_13432_ _13431_/X rdata[30] _13516_/S VGND VGND VPWR VPWR _13432_/X sky130_fd_sc_hd__mux2_1
X_10644_ _14760_/Q _10637_/X _10415_/X _10638_/X VGND VGND VPWR VPWR _14760_/D sky130_fd_sc_hd__a22o_1
XFILLER_10_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13363_ _13364_/X _12519_/B _13415_/S VGND VGND VPWR VPWR _13363_/X sky130_fd_sc_hd__mux2_1
X_10575_ _10584_/A VGND VGND VPWR VPWR _10575_/X sky130_fd_sc_hd__buf_1
X_15102_ _09316_/X _15102_/D VGND VGND VPWR VPWR _15102_/Q sky130_fd_sc_hd__dfxtp_1
X_12314_ _12432_/D _12431_/A _12745_/A _12357_/B VGND VGND VPWR VPWR _12342_/B sky130_fd_sc_hd__a211oi_4
X_13294_ _13335_/X _13333_/X _13408_/S VGND VGND VPWR VPWR _13294_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15033_ _09576_/X _15033_/D VGND VGND VPWR VPWR _15033_/Q sky130_fd_sc_hd__dfxtp_1
X_12245_ _12243_/X _12081_/A _12825_/A _12130_/A VGND VGND VPWR VPWR _12246_/B sky130_fd_sc_hd__o22a_1
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12176_ _12725_/A _12271_/B _12175_/Y VGND VGND VPWR VPWR _12684_/A sky130_fd_sc_hd__a21oi_2
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11127_ _14645_/Q _11120_/X _11126_/X _11123_/X VGND VGND VPWR VPWR _14645_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11058_ _11070_/A VGND VGND VPWR VPWR _11058_/X sky130_fd_sc_hd__clkbuf_1
X_10009_ _14929_/Q _09998_/X _10008_/X _10000_/X VGND VGND VPWR VPWR _14929_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14817_ _10445_/X _14817_/D VGND VGND VPWR VPWR _14817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_opt_1_clk _14315_/CLK VGND VGND VPWR VPWR _14375_/CLK sky130_fd_sc_hd__clkbuf_16
X_14748_ _10700_/X _14748_/D VGND VGND VPWR VPWR _14748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14679_ _10991_/X _14679_/D VGND VGND VPWR VPWR _14679_/Q sky130_fd_sc_hd__dfxtp_1
X_07220_ _07220_/A VGND VGND VPWR VPWR _07220_/Y sky130_fd_sc_hd__inv_2
X_07151_ _13091_/X VGND VGND VPWR VPWR _07237_/A sky130_fd_sc_hd__inv_2
XFILLER_105_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07984_ _07984_/A VGND VGND VPWR VPWR _07984_/X sky130_fd_sc_hd__buf_1
X_09723_ _15005_/Q _09715_/X _09559_/X _09718_/X VGND VGND VPWR VPWR _15005_/D sky130_fd_sc_hd__a22o_1
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09654_ _09684_/A VGND VGND VPWR VPWR _09665_/A sky130_fd_sc_hd__buf_1
XFILLER_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08605_ _08605_/A VGND VGND VPWR VPWR _08612_/A sky130_fd_sc_hd__buf_1
XFILLER_82_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09585_ _15032_/Q _09577_/X _09584_/X _09580_/X VGND VGND VPWR VPWR _15032_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08536_ _15301_/Q _08520_/X _08535_/X _08524_/X VGND VGND VPWR VPWR _15301_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08467_ _08467_/A VGND VGND VPWR VPWR _08467_/X sky130_fd_sc_hd__buf_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07418_ _07419_/A _13587_/X VGND VGND VPWR VPWR _15577_/D sky130_fd_sc_hd__and2_1
X_08398_ _08416_/A VGND VGND VPWR VPWR _08411_/A sky130_fd_sc_hd__buf_1
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07349_ _07353_/A _07349_/B VGND VGND VPWR VPWR _15599_/D sky130_fd_sc_hd__nor2_1
XFILLER_149_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10360_ _14837_/Q _10353_/X _10359_/X _10356_/X VGND VGND VPWR VPWR _14837_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09019_ _09021_/A VGND VGND VPWR VPWR _09019_/X sky130_fd_sc_hd__clkbuf_1
X_10291_ _10302_/A VGND VGND VPWR VPWR _10291_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12030_ _12040_/A _12037_/A _12030_/C _12040_/B VGND VGND VPWR VPWR _12031_/A sky130_fd_sc_hd__or4_4
XFILLER_88_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13981_ _13977_/X _13978_/X _13979_/X _13980_/X _14397_/Q _14398_/Q VGND VGND VPWR
+ VPWR _13981_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12932_ _12828_/X _12825_/X _12924_/C _12931_/X VGND VGND VPWR VPWR _12933_/B sky130_fd_sc_hd__o22a_1
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15651_ _15652_/CLK _15651_/D VGND VGND VPWR VPWR _15651_/Q sky130_fd_sc_hd__dfxtp_1
X_12863_ _12863_/A VGND VGND VPWR VPWR _12863_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14602_ _11293_/X _14602_/D VGND VGND VPWR VPWR _14602_/Q sky130_fd_sc_hd__dfxtp_1
X_11814_ _11814_/A VGND VGND VPWR VPWR _11876_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15582_ _15591_/CLK _15582_/D VGND VGND VPWR VPWR _15582_/Q sky130_fd_sc_hd__dfxtp_1
X_12794_ _12747_/Y _12201_/A _12686_/X _12209_/B _12681_/X VGND VGND VPWR VPWR _12794_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14533_ _11563_/X _14533_/D VGND VGND VPWR VPWR _14533_/Q sky130_fd_sc_hd__dfxtp_1
X_11745_ _14483_/Q _11743_/X _11502_/X _11744_/X VGND VGND VPWR VPWR _14483_/D sky130_fd_sc_hd__a22o_1
X_14464_ _11808_/X _14464_/D VGND VGND VPWR VPWR _14464_/Q sky130_fd_sc_hd__dfxtp_1
X_11676_ _11678_/A VGND VGND VPWR VPWR _11676_/X sky130_fd_sc_hd__clkbuf_1
X_13415_ _13417_/X _13416_/X _13415_/S VGND VGND VPWR VPWR _13415_/X sky130_fd_sc_hd__mux2_1
X_10627_ _10646_/A VGND VGND VPWR VPWR _10627_/X sky130_fd_sc_hd__buf_1
X_14395_ _14395_/CLK instruction[20] VGND VGND VPWR VPWR _14395_/Q sky130_fd_sc_hd__dfxtp_4
X_13346_ _13399_/X _13397_/X _13415_/S VGND VGND VPWR VPWR _13346_/X sky130_fd_sc_hd__mux2_1
X_10558_ _14785_/Q _10550_/X _10303_/X _10553_/X VGND VGND VPWR VPWR _14785_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13277_ _12785_/A _12775_/X _15561_/Q VGND VGND VPWR VPWR _13277_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10489_ _14805_/Q _10484_/X _10359_/X _10486_/X VGND VGND VPWR VPWR _14805_/D sky130_fd_sc_hd__a22o_1
X_15016_ _09670_/X _15016_/D VGND VGND VPWR VPWR _15016_/Q sky130_fd_sc_hd__dfxtp_1
X_12228_ _12228_/A VGND VGND VPWR VPWR _12228_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12159_ _12155_/X _12157_/X _12708_/A _12148_/X VGND VGND VPWR VPWR _12160_/B sky130_fd_sc_hd__o22a_1
XFILLER_111_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09370_ _09370_/A VGND VGND VPWR VPWR _09370_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08321_ _15337_/Q _08316_/X _08069_/X _08317_/X VGND VGND VPWR VPWR _15337_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08252_ _08261_/A VGND VGND VPWR VPWR _08252_/X sky130_fd_sc_hd__buf_1
XFILLER_138_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07203_ _13112_/X _07202_/Y _07198_/X _07173_/B VGND VGND VPWR VPWR _15658_/D sky130_fd_sc_hd__o211a_1
X_08183_ _08204_/A VGND VGND VPWR VPWR _08183_/X sky130_fd_sc_hd__buf_1
XFILLER_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07134_ _13110_/X VGND VGND VPWR VPWR _07264_/B sky130_fd_sc_hd__inv_2
XFILLER_106_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07967_ _14329_/Q VGND VGND VPWR VPWR _07968_/A sky130_fd_sc_hd__buf_1
XFILLER_68_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09706_ _15010_/Q _09702_/X _09527_/X _09705_/X VGND VGND VPWR VPWR _15010_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07898_ _07897_/A _07897_/B _07893_/X _07897_/Y VGND VGND VPWR VPWR _15432_/D sky130_fd_sc_hd__o211a_1
X_09637_ _10389_/A VGND VGND VPWR VPWR _09637_/X sky130_fd_sc_hd__buf_1
XFILLER_55_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09568_ _10707_/A VGND VGND VPWR VPWR _10332_/A sky130_fd_sc_hd__buf_1
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ _08526_/A VGND VGND VPWR VPWR _08519_/X sky130_fd_sc_hd__clkbuf_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09499_ _09499_/A VGND VGND VPWR VPWR _09504_/A sky130_fd_sc_hd__buf_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11530_ _11554_/A VGND VGND VPWR VPWR _11530_/X sky130_fd_sc_hd__buf_1
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11461_ _11466_/A VGND VGND VPWR VPWR _11461_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13200_ _13201_/X _13221_/X _13408_/S VGND VGND VPWR VPWR _13200_/X sky130_fd_sc_hd__mux2_1
X_10412_ _14825_/Q _10406_/X _10411_/X _10408_/X VGND VGND VPWR VPWR _14825_/D sky130_fd_sc_hd__a22o_1
X_14180_ _14958_/Q _15054_/Q _15022_/Q _15086_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14180_/X sky130_fd_sc_hd__mux4_2
X_11392_ _11392_/A VGND VGND VPWR VPWR _11392_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13131_ _12610_/X _13016_/Y _13152_/S VGND VGND VPWR VPWR _13131_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10343_ _10343_/A VGND VGND VPWR VPWR _10343_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13062_ _12872_/Y _15564_/Q _13090_/S VGND VGND VPWR VPWR _13062_/X sky130_fd_sc_hd__mux2_1
X_10274_ _10290_/A VGND VGND VPWR VPWR _10279_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12013_ _12017_/A VGND VGND VPWR VPWR _12013_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13964_ _15171_/Q _15139_/Q _14755_/Q _14787_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13964_/X sky130_fd_sc_hd__mux4_1
X_12915_ _12778_/X _12204_/X _12773_/A _12779_/A VGND VGND VPWR VPWR _12919_/A sky130_fd_sc_hd__o22a_1
XFILLER_34_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13895_ _15114_/Q _15338_/Q _15306_/Q _15274_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13895_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15634_ _15666_/CLK _15634_/D VGND VGND VPWR VPWR pc[29] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12846_ _12846_/A _12846_/B VGND VGND VPWR VPWR _12846_/X sky130_fd_sc_hd__or2_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15565_ _15566_/CLK _15565_/D VGND VGND VPWR VPWR _15565_/Q sky130_fd_sc_hd__dfxtp_4
X_12777_ _12746_/X _12776_/X _12746_/X _12776_/X VGND VGND VPWR VPWR _12777_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14516_ _11628_/X _14516_/D VGND VGND VPWR VPWR _14516_/Q sky130_fd_sc_hd__dfxtp_1
X_11728_ _14488_/Q _11722_/X _11479_/X _11723_/X VGND VGND VPWR VPWR _14488_/D sky130_fd_sc_hd__a22o_1
X_15496_ _15591_/CLK _15496_/D VGND VGND VPWR VPWR wdata[22] sky130_fd_sc_hd__dfxtp_4
XFILLER_147_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14447_ _11868_/X _14447_/D VGND VGND VPWR VPWR _14447_/Q sky130_fd_sc_hd__dfxtp_1
X_11659_ _14507_/Q _11652_/X _11537_/X _11654_/X VGND VGND VPWR VPWR _14507_/D sky130_fd_sc_hd__a22o_1
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14378_ _14391_/CLK instruction[7] VGND VGND VPWR VPWR _14378_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13329_ _13330_/X _12520_/B _13408_/S VGND VGND VPWR VPWR _13329_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08870_ _15215_/Q _08864_/X _08869_/X _08866_/X VGND VGND VPWR VPWR _15215_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07821_ _07821_/A _07779_/A VGND VGND VPWR VPWR _07822_/A sky130_fd_sc_hd__or2b_1
XFILLER_57_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07752_ _07895_/B VGND VGND VPWR VPWR _07752_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07683_ _13134_/X VGND VGND VPWR VPWR _07683_/X sky130_fd_sc_hd__buf_1
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09422_ _09422_/A VGND VGND VPWR VPWR _09422_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09353_ _09383_/A VGND VGND VPWR VPWR _09372_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_33_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08304_ _08304_/A VGND VGND VPWR VPWR _08304_/X sky130_fd_sc_hd__clkbuf_1
X_09284_ _09284_/A VGND VGND VPWR VPWR _09284_/X sky130_fd_sc_hd__buf_1
XFILLER_21_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08235_ _15361_/Q _08227_/X _07936_/X _08230_/X VGND VGND VPWR VPWR _15361_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08166_ _15379_/Q _08164_/X _08016_/X _08165_/X VGND VGND VPWR VPWR _15379_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07117_ _15513_/Q VGND VGND VPWR VPWR _12040_/A sky130_fd_sc_hd__buf_1
XFILLER_107_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08097_ _08097_/A VGND VGND VPWR VPWR _08097_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08999_ _15182_/Q _08993_/X _08873_/X _08994_/X VGND VGND VPWR VPWR _15182_/D sky130_fd_sc_hd__a22o_1
XFILLER_75_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10961_ _10961_/A VGND VGND VPWR VPWR _10961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12700_ _12783_/A VGND VGND VPWR VPWR _12706_/A sky130_fd_sc_hd__buf_1
XFILLER_16_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13680_ _14976_/Q _15072_/Q _15040_/Q _15104_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13680_/X sky130_fd_sc_hd__mux4_2
X_10892_ _10892_/A VGND VGND VPWR VPWR _10899_/A sky130_fd_sc_hd__buf_1
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12631_ _12611_/X _12946_/B _12600_/X _13214_/X _12451_/X VGND VGND VPWR VPWR _12632_/B
+ sky130_fd_sc_hd__o32a_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ _08270_/X _15350_/D VGND VGND VPWR VPWR _15350_/Q sky130_fd_sc_hd__dfxtp_1
X_12562_ _12546_/A _12561_/Y _12553_/A VGND VGND VPWR VPWR wstrobe[3] sky130_fd_sc_hd__o21a_2
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14301_ _15469_/CLK _15468_/Q VGND VGND VPWR VPWR _14301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11513_ _11513_/A VGND VGND VPWR VPWR _11513_/X sky130_fd_sc_hd__buf_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15281_ _08612_/X _15281_/D VGND VGND VPWR VPWR _15281_/Q sky130_fd_sc_hd__dfxtp_1
X_12493_ _12493_/A VGND VGND VPWR VPWR _12493_/X sky130_fd_sc_hd__clkbuf_4
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ _15208_/Q _14536_/Q _14984_/Q _15400_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14232_/X sky130_fd_sc_hd__mux4_2
X_11444_ _14560_/Q _11430_/X _11443_/X _11434_/X VGND VGND VPWR VPWR _14560_/D sky130_fd_sc_hd__a22o_1
X_14163_ _14671_/Q _15247_/Q _14735_/Q _14703_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14163_/X sky130_fd_sc_hd__mux4_2
X_11375_ _11385_/A VGND VGND VPWR VPWR _11375_/X sky130_fd_sc_hd__buf_1
X_13114_ _15660_/Q data_address[25] _15667_/Q VGND VGND VPWR VPWR _13114_/X sky130_fd_sc_hd__mux2_1
X_10326_ _10331_/A VGND VGND VPWR VPWR _10326_/X sky130_fd_sc_hd__clkbuf_1
X_14094_ _15190_/Q _15158_/Q _14774_/Q _14806_/Q _14238_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14094_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13045_ wdata[18] rdata[18] _13058_/S VGND VGND VPWR VPWR _14322_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10257_ _10280_/A VGND VGND VPWR VPWR _10257_/X sky130_fd_sc_hd__buf_1
XFILLER_67_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10188_ _10201_/A VGND VGND VPWR VPWR _10193_/A sky130_fd_sc_hd__buf_1
XFILLER_79_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14996_ _09752_/X _14996_/D VGND VGND VPWR VPWR _14996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13947_ _14629_/Q _14597_/Q _14565_/Q _15365_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13947_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13878_ _14508_/Q _14476_/Q _14444_/Q _14412_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13878_/X sky130_fd_sc_hd__mux4_2
XFILLER_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15617_ _15647_/CLK _15617_/D VGND VGND VPWR VPWR pc[12] sky130_fd_sc_hd__dfxtp_1
X_12829_ _12829_/A VGND VGND VPWR VPWR _12829_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15548_ _15579_/CLK _15548_/D VGND VGND VPWR VPWR _15548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15479_ _15566_/CLK _15479_/D VGND VGND VPWR VPWR wdata[5] sky130_fd_sc_hd__dfxtp_4
X_08020_ _14319_/Q VGND VGND VPWR VPWR _08021_/A sky130_fd_sc_hd__buf_1
XFILLER_144_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09971_ _09976_/A VGND VGND VPWR VPWR _09971_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08922_ _08936_/A VGND VGND VPWR VPWR _08922_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08853_ _08866_/A VGND VGND VPWR VPWR _08853_/X sky130_fd_sc_hd__buf_1
XFILLER_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07804_ _07804_/A _07804_/B VGND VGND VPWR VPWR _07805_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08784_ _08796_/A VGND VGND VPWR VPWR _08800_/A sky130_fd_sc_hd__inv_2
XFILLER_85_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07735_ _13143_/X _07728_/B _07728_/Y VGND VGND VPWR VPWR _07874_/A sky130_fd_sc_hd__a21oi_1
XFILLER_65_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07666_ _07798_/B VGND VGND VPWR VPWR _07666_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09405_ _09407_/A VGND VGND VPWR VPWR _09405_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07597_ _07599_/A _13070_/X VGND VGND VPWR VPWR _15485_/D sky130_fd_sc_hd__and2_1
X_09336_ _09336_/A VGND VGND VPWR VPWR _09336_/X sky130_fd_sc_hd__buf_1
XFILLER_138_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09267_ _09267_/A VGND VGND VPWR VPWR _09267_/X sky130_fd_sc_hd__buf_1
XFILLER_138_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08218_ _09923_/B VGND VGND VPWR VPWR _09294_/B sky130_fd_sc_hd__clkbuf_1
X_09198_ _15129_/Q _09195_/X _09196_/X _09197_/X VGND VGND VPWR VPWR _15129_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08149_ _15383_/Q _08143_/X _07994_/X _08144_/X VGND VGND VPWR VPWR _15383_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11160_ _11186_/A VGND VGND VPWR VPWR _11160_/X sky130_fd_sc_hd__buf_1
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10111_ _10111_/A VGND VGND VPWR VPWR _10111_/X sky130_fd_sc_hd__clkbuf_1
X_11091_ _11459_/A VGND VGND VPWR VPWR _11091_/X sky130_fd_sc_hd__buf_1
XFILLER_96_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10042_ _10411_/A VGND VGND VPWR VPWR _10042_/X sky130_fd_sc_hd__buf_1
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14850_ _10293_/X _14850_/D VGND VGND VPWR VPWR _14850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13801_ _13797_/X _13798_/X _13799_/X _13800_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13801_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14781_ _10572_/X _14781_/D VGND VGND VPWR VPWR _14781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11993_ _14411_/Q _11986_/X _08059_/A _11988_/X VGND VGND VPWR VPWR _14411_/D sky130_fd_sc_hd__a22o_1
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13732_ _15226_/Q _14554_/Q _15002_/Q _15418_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13732_/X sky130_fd_sc_hd__mux4_1
X_10944_ _10948_/A VGND VGND VPWR VPWR _10944_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13663_ _14689_/Q _15265_/Q _14753_/Q _14721_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13663_/X sky130_fd_sc_hd__mux4_2
X_10875_ _10875_/A VGND VGND VPWR VPWR _10875_/X sky130_fd_sc_hd__buf_1
XFILLER_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15402_ _08061_/X _15402_/D VGND VGND VPWR VPWR _15402_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12614_ _12579_/X _12613_/X _12579_/X _12613_/X VGND VGND VPWR VPWR _12614_/Y sky130_fd_sc_hd__a2bb2oi_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13594_ _13593_/X _14318_/D _15506_/Q VGND VGND VPWR VPWR _13594_/X sky130_fd_sc_hd__mux2_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15333_ _08332_/X _15333_/D VGND VGND VPWR VPWR _15333_/Q sky130_fd_sc_hd__dfxtp_1
X_12545_ _12545_/A _12551_/A _12545_/C VGND VGND VPWR VPWR _12546_/A sky130_fd_sc_hd__and3_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15264_ _08674_/X _15264_/D VGND VGND VPWR VPWR _15264_/Q sky130_fd_sc_hd__dfxtp_1
X_12476_ _12480_/A _12480_/B _12475_/X VGND VGND VPWR VPWR _12476_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14215_ _15114_/Q _15338_/Q _15306_/Q _15274_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14215_/X sky130_fd_sc_hd__mux4_1
XANTENNA_5 data_address[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11427_ _11436_/A VGND VGND VPWR VPWR _11427_/X sky130_fd_sc_hd__clkbuf_1
X_15195_ _08957_/X _15195_/D VGND VGND VPWR VPWR _15195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14146_ _14142_/X _14143_/X _14144_/X _14145_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14146_/X sky130_fd_sc_hd__mux4_2
X_11358_ _11362_/A VGND VGND VPWR VPWR _11358_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10309_ _14848_/Q _10296_/X _10308_/X _10300_/X VGND VGND VPWR VPWR _14848_/D sky130_fd_sc_hd__a22o_1
X_14077_ _14648_/Q _14616_/Q _14584_/Q _15384_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14077_/X sky130_fd_sc_hd__mux4_2
X_11289_ _14604_/Q _11284_/X _11166_/X _11286_/X VGND VGND VPWR VPWR _14604_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13028_ wdata[1] rdata[1] _13058_/S VGND VGND VPWR VPWR _14305_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14979_ _09807_/X _14979_/D VGND VGND VPWR VPWR _14979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07520_ _07635_/A _14372_/Q VGND VGND VPWR VPWR _15508_/D sky130_fd_sc_hd__or2_1
XFILLER_35_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07451_ _07451_/A _13445_/X VGND VGND VPWR VPWR _15555_/D sky130_fd_sc_hd__and2_1
XFILLER_50_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07382_ _07385_/B VGND VGND VPWR VPWR _07382_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09121_ _09125_/A VGND VGND VPWR VPWR _09121_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09052_ _09052_/A VGND VGND VPWR VPWR _09115_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08003_ _15414_/Q _07998_/X _08000_/X _08002_/X VGND VGND VPWR VPWR _15414_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09954_ _10324_/A VGND VGND VPWR VPWR _09954_/X sky130_fd_sc_hd__buf_1
X_08905_ _09275_/A VGND VGND VPWR VPWR _08905_/X sky130_fd_sc_hd__buf_1
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09885_ _09885_/A VGND VGND VPWR VPWR _09885_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08836_ _08843_/A VGND VGND VPWR VPWR _08836_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08767_ _15238_/Q _08762_/X _08529_/X _08763_/X VGND VGND VPWR VPWR _15238_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07718_ _07871_/B _07868_/A VGND VGND VPWR VPWR _07774_/C sky130_fd_sc_hd__or2_1
X_08698_ _15259_/Q _08693_/X _08396_/X _08694_/X VGND VGND VPWR VPWR _15259_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07649_ _07701_/A VGND VGND VPWR VPWR _07650_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10660_ _10670_/A VGND VGND VPWR VPWR _10660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09319_ _15101_/Q _09311_/X _09180_/X _09314_/X VGND VGND VPWR VPWR _15101_/D sky130_fd_sc_hd__a22o_1
X_10591_ _10595_/A VGND VGND VPWR VPWR _10591_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12330_ _12330_/A VGND VGND VPWR VPWR _12330_/X sky130_fd_sc_hd__buf_1
XFILLER_108_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12261_ _12261_/A VGND VGND VPWR VPWR _12261_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14000_ _14976_/Q _15072_/Q _15040_/Q _15104_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _14000_/X sky130_fd_sc_hd__mux4_2
XFILLER_123_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11212_ _11214_/A VGND VGND VPWR VPWR _11212_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12192_ _12762_/A _12190_/B _12191_/Y VGND VGND VPWR VPWR _12749_/A sky130_fd_sc_hd__a21oi_4
XFILLER_150_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11143_ _11151_/A VGND VGND VPWR VPWR _11143_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11074_ _11086_/A VGND VGND VPWR VPWR _11074_/X sky130_fd_sc_hd__clkbuf_1
X_14902_ _10115_/X _14902_/D VGND VGND VPWR VPWR _14902_/Q sky130_fd_sc_hd__dfxtp_1
X_10025_ _10394_/A VGND VGND VPWR VPWR _10025_/X sky130_fd_sc_hd__buf_1
XFILLER_49_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14833_ _10374_/X _14833_/D VGND VGND VPWR VPWR _14833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14764_ _10632_/X _14764_/D VGND VGND VPWR VPWR _14764_/Q sky130_fd_sc_hd__dfxtp_1
X_11976_ _11976_/A VGND VGND VPWR VPWR _11976_/X sky130_fd_sc_hd__buf_1
XFILLER_91_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13715_ _15132_/Q _15356_/Q _15324_/Q _15292_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13715_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10927_ _10929_/A VGND VGND VPWR VPWR _10927_/X sky130_fd_sc_hd__clkbuf_1
X_14695_ _10935_/X _14695_/D VGND VGND VPWR VPWR _14695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13646_ _13645_/X _14305_/D _15506_/Q VGND VGND VPWR VPWR _13646_/X sky130_fd_sc_hd__mux2_1
X_10858_ _10860_/A VGND VGND VPWR VPWR _10858_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13577_ _13576_/X _13581_/A1 _13649_/S VGND VGND VPWR VPWR _13577_/X sky130_fd_sc_hd__mux2_1
X_10789_ _14732_/Q _10780_/X _10788_/X _10784_/X VGND VGND VPWR VPWR _14732_/D sky130_fd_sc_hd__a22o_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15316_ _08439_/X _15316_/D VGND VGND VPWR VPWR _15316_/Q sky130_fd_sc_hd__dfxtp_1
X_12528_ _15592_/Q _12962_/B _12501_/X _12527_/X VGND VGND VPWR VPWR _12528_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15247_ _08736_/X _15247_/D VGND VGND VPWR VPWR _15247_/Q sky130_fd_sc_hd__dfxtp_1
X_12459_ _12846_/B _12459_/B VGND VGND VPWR VPWR _12459_/X sky130_fd_sc_hd__or2_1
XFILLER_99_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15178_ _09015_/X _15178_/D VGND VGND VPWR VPWR _15178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14129_ _14835_/Q _14867_/Q _14899_/Q _14931_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14129_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09670_ _09680_/A VGND VGND VPWR VPWR _09670_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08621_ _15279_/Q _08617_/X _08472_/X _08618_/X VGND VGND VPWR VPWR _15279_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08552_ _08552_/A VGND VGND VPWR VPWR _08552_/X sky130_fd_sc_hd__buf_1
X_07503_ _14384_/Q VGND VGND VPWR VPWR _12563_/A sky130_fd_sc_hd__inv_2
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08483_ _14314_/Q VGND VGND VPWR VPWR _10781_/A sky130_fd_sc_hd__buf_1
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07434_ _07460_/A VGND VGND VPWR VPWR _07443_/A sky130_fd_sc_hd__buf_1
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07365_ _14398_/Q VGND VGND VPWR VPWR _07366_/A sky130_fd_sc_hd__inv_2
X_09104_ _15153_/Q _09095_/X _08861_/X _09096_/X VGND VGND VPWR VPWR _15153_/D sky130_fd_sc_hd__a22o_1
X_07296_ _07559_/C _14376_/Q _07559_/A _07559_/B VGND VGND VPWR VPWR _07297_/A sky130_fd_sc_hd__or4_4
X_09035_ _15172_/Q _08929_/A _08916_/X _08932_/A VGND VGND VPWR VPWR _15172_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09937_ _09949_/A VGND VGND VPWR VPWR _09937_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09868_ _09877_/A VGND VGND VPWR VPWR _09868_/X sky130_fd_sc_hd__buf_1
XFILLER_133_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08819_ _08858_/A VGND VGND VPWR VPWR _08846_/A sky130_fd_sc_hd__buf_2
XFILLER_46_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09799_ _14983_/Q _09797_/X _09677_/X _09798_/X VGND VGND VPWR VPWR _14983_/D sky130_fd_sc_hd__a22o_1
XFILLER_133_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_203 _13570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11830_ _11839_/A VGND VGND VPWR VPWR _11837_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_214 _13776_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_225 _08431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_236 _10790_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_247 _11895_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_258 _15538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11761_ _14478_/Q _11752_/X _11523_/X _11753_/X VGND VGND VPWR VPWR _14478_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13500_ _13896_/X _13901_/X _13521_/S VGND VGND VPWR VPWR _13500_/X sky130_fd_sc_hd__mux2_1
X_10712_ _10712_/A VGND VGND VPWR VPWR _11471_/A sky130_fd_sc_hd__buf_1
X_14480_ _11751_/X _14480_/D VGND VGND VPWR VPWR _14480_/Q sky130_fd_sc_hd__dfxtp_1
X_11692_ _14498_/Q _11688_/X _11431_/X _11691_/X VGND VGND VPWR VPWR _14498_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13431_ _13666_/X _13671_/X _13521_/S VGND VGND VPWR VPWR _13431_/X sky130_fd_sc_hd__mux2_1
X_10643_ _10645_/A VGND VGND VPWR VPWR _10643_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13362_ _13365_/X _13363_/X _13408_/S VGND VGND VPWR VPWR _13362_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10574_ _10574_/A VGND VGND VPWR VPWR _10574_/X sky130_fd_sc_hd__clkbuf_1
X_15101_ _09318_/X _15101_/D VGND VGND VPWR VPWR _15101_/Q sky130_fd_sc_hd__dfxtp_1
X_12313_ _12432_/D _12431_/A VGND VGND VPWR VPWR _12357_/B sky130_fd_sc_hd__nor2_2
X_13293_ _13332_/X _13330_/X _13408_/S VGND VGND VPWR VPWR _13293_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15032_ _09582_/X _15032_/D VGND VGND VPWR VPWR _15032_/Q sky130_fd_sc_hd__dfxtp_1
X_12244_ _15567_/Q VGND VGND VPWR VPWR _12825_/A sky130_fd_sc_hd__inv_2
XFILLER_108_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12175_ _12271_/A _12271_/B VGND VGND VPWR VPWR _12175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11126_ _11494_/A VGND VGND VPWR VPWR _11126_/X sky130_fd_sc_hd__buf_1
XFILLER_122_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11057_ _11089_/A VGND VGND VPWR VPWR _11070_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10008_ _10375_/A VGND VGND VPWR VPWR _10008_/X sky130_fd_sc_hd__buf_1
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14816_ _10447_/X _14816_/D VGND VGND VPWR VPWR _14816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14747_ _10706_/X _14747_/D VGND VGND VPWR VPWR _14747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11959_ _14422_/Q _11956_/X _08000_/A _11958_/X VGND VGND VPWR VPWR _14422_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14678_ _10993_/X _14678_/D VGND VGND VPWR VPWR _14678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13629_ _13628_/X _07352_/Y _13641_/S VGND VGND VPWR VPWR _13629_/X sky130_fd_sc_hd__mux2_1
Xrepeater50 _14060_/S0 VGND VGND VPWR VPWR _07387_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_20_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07150_ _13092_/X VGND VGND VPWR VPWR _07236_/A sky130_fd_sc_hd__inv_2
XFILLER_9_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07983_ _07983_/A VGND VGND VPWR VPWR _07983_/X sky130_fd_sc_hd__buf_1
XFILLER_101_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09722_ _09722_/A VGND VGND VPWR VPWR _09722_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09653_ _09733_/A VGND VGND VPWR VPWR _09684_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08604_ _15284_/Q _08597_/X _08442_/X _08599_/X VGND VGND VPWR VPWR _15284_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09584_ _10344_/A VGND VGND VPWR VPWR _09584_/X sky130_fd_sc_hd__buf_1
XFILLER_36_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08535_ _09284_/A VGND VGND VPWR VPWR _08535_/X sky130_fd_sc_hd__buf_1
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08466_ _09236_/A VGND VGND VPWR VPWR _08466_/X sky130_fd_sc_hd__buf_1
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ _07419_/A _13583_/X VGND VGND VPWR VPWR _15578_/D sky130_fd_sc_hd__and2_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08397_ _15323_/Q _08387_/X _08396_/X _08391_/X VGND VGND VPWR VPWR _15323_/D sky130_fd_sc_hd__a22o_1
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07348_ _07349_/B VGND VGND VPWR VPWR _07348_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07279_ _07283_/A VGND VGND VPWR VPWR _07282_/A sky130_fd_sc_hd__buf_1
X_09018_ _15178_/Q _09016_/X _08891_/X _09017_/X VGND VGND VPWR VPWR _15178_/D sky130_fd_sc_hd__a22o_1
X_10290_ _10290_/A VGND VGND VPWR VPWR _10302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13980_ _14978_/Q _15074_/Q _15042_/Q _15106_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13980_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12931_ _12852_/A _12854_/X _12924_/A _12842_/X _12847_/B VGND VGND VPWR VPWR _12931_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15650_ _15652_/CLK _15650_/D VGND VGND VPWR VPWR _15650_/Q sky130_fd_sc_hd__dfxtp_1
X_12862_ _12862_/A VGND VGND VPWR VPWR _12875_/B sky130_fd_sc_hd__buf_2
XFILLER_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11813_ _11834_/A VGND VGND VPWR VPWR _11813_/X sky130_fd_sc_hd__buf_1
X_14601_ _11297_/X _14601_/D VGND VGND VPWR VPWR _14601_/Q sky130_fd_sc_hd__dfxtp_1
X_15581_ _15592_/CLK _15581_/D VGND VGND VPWR VPWR _15581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12793_ _12791_/X _12195_/X _12713_/X _12792_/X VGND VGND VPWR VPWR _12793_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_42_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14532_ _11566_/X _14532_/D VGND VGND VPWR VPWR _14532_/Q sky130_fd_sc_hd__dfxtp_1
X_11744_ _11753_/A VGND VGND VPWR VPWR _11744_/X sky130_fd_sc_hd__buf_1
XFILLER_14_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14463_ _11810_/X _14463_/D VGND VGND VPWR VPWR _14463_/Q sky130_fd_sc_hd__dfxtp_1
X_11675_ _14503_/Q _11673_/X _11553_/X _11674_/X VGND VGND VPWR VPWR _14503_/D sky130_fd_sc_hd__a22o_1
XFILLER_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13414_ _12775_/X _12785_/A _13418_/S VGND VGND VPWR VPWR _13414_/X sky130_fd_sc_hd__mux2_1
X_10626_ _10626_/A VGND VGND VPWR VPWR _10646_/A sky130_fd_sc_hd__clkbuf_2
X_14394_ _14399_/CLK instruction[31] VGND VGND VPWR VPWR _14394_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13345_ _13346_/X _12488_/B _13408_/S VGND VGND VPWR VPWR _13345_/X sky130_fd_sc_hd__mux2_1
X_10557_ _10561_/A VGND VGND VPWR VPWR _10557_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13276_ _13277_/X _13288_/X _15562_/Q VGND VGND VPWR VPWR _13276_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10488_ _10490_/A VGND VGND VPWR VPWR _10488_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15015_ _09674_/X _15015_/D VGND VGND VPWR VPWR _15015_/Q sky130_fd_sc_hd__dfxtp_1
X_12227_ _12885_/A _12225_/X _13354_/X _12892_/A VGND VGND VPWR VPWR _12228_/A sky130_fd_sc_hd__o22a_1
XFILLER_142_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12158_ _15575_/Q VGND VGND VPWR VPWR _12708_/A sky130_fd_sc_hd__inv_2
XFILLER_78_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11109_ _11109_/A VGND VGND VPWR VPWR _11109_/X sky130_fd_sc_hd__buf_1
X_12089_ _12598_/A _12585_/A VGND VGND VPWR VPWR _12089_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08320_ _08324_/A VGND VGND VPWR VPWR _08320_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08251_ _08251_/A VGND VGND VPWR VPWR _08251_/X sky130_fd_sc_hd__clkbuf_1
X_07202_ _07202_/A VGND VGND VPWR VPWR _07202_/Y sky130_fd_sc_hd__inv_2
X_08182_ _08182_/A VGND VGND VPWR VPWR _08204_/A sky130_fd_sc_hd__clkbuf_2
X_07133_ _13111_/X VGND VGND VPWR VPWR _07263_/B sky130_fd_sc_hd__inv_2
XFILLER_106_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07966_ _07981_/A VGND VGND VPWR VPWR _07966_/X sky130_fd_sc_hd__buf_1
XFILLER_75_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09705_ _09705_/A VGND VGND VPWR VPWR _09705_/X sky130_fd_sc_hd__buf_1
XFILLER_28_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07897_ _07897_/A _07897_/B VGND VGND VPWR VPWR _07897_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09636_ _10775_/A VGND VGND VPWR VPWR _10389_/A sky130_fd_sc_hd__buf_1
XFILLER_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09567_ _09567_/A VGND VGND VPWR VPWR _09567_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08518_ _15304_/Q _08502_/X _08517_/X _08506_/X VGND VGND VPWR VPWR _15304_/D sky130_fd_sc_hd__a22o_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09498_ _15050_/Q _09496_/X _09263_/X _09497_/X VGND VGND VPWR VPWR _15050_/D sky130_fd_sc_hd__a22o_1
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08449_ _08467_/A VGND VGND VPWR VPWR _08449_/X sky130_fd_sc_hd__buf_1
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11460_ _14557_/Q _11448_/X _11459_/X _11452_/X VGND VGND VPWR VPWR _14557_/D sky130_fd_sc_hd__a22o_1
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10411_ _10411_/A VGND VGND VPWR VPWR _10411_/X sky130_fd_sc_hd__buf_1
X_11391_ _14574_/Q _11384_/X _11156_/X _11385_/X VGND VGND VPWR VPWR _14574_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13130_ _12577_/X _13017_/Y _13152_/S VGND VGND VPWR VPWR _13130_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10342_ _14841_/Q _10339_/X _10340_/X _10341_/X VGND VGND VPWR VPWR _14841_/D sky130_fd_sc_hd__a22o_1
XFILLER_125_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13061_ _12881_/Y _15563_/Q _13076_/S VGND VGND VPWR VPWR _13061_/X sky130_fd_sc_hd__mux2_2
XFILLER_124_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10273_ _10346_/A VGND VGND VPWR VPWR _10290_/A sky130_fd_sc_hd__buf_1
XFILLER_79_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12012_ _12012_/A VGND VGND VPWR VPWR _12017_/A sky130_fd_sc_hd__buf_1
XFILLER_78_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13963_ _14659_/Q _15235_/Q _14723_/Q _14691_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13963_/X sky130_fd_sc_hd__mux4_2
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12914_ _12941_/A _12914_/B _12914_/C _12913_/X VGND VGND VPWR VPWR _12957_/D sky130_fd_sc_hd__or4b_4
XFILLER_74_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13894_ _15178_/Q _15146_/Q _14762_/Q _14794_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13894_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15633_ _15666_/CLK _15633_/D VGND VGND VPWR VPWR pc[28] sky130_fd_sc_hd__dfxtp_2
XFILLER_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12845_ _12842_/X _12251_/X _12501_/X _12844_/X VGND VGND VPWR VPWR _12845_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_61_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12776_ _12775_/A _12199_/A _12686_/X _12209_/B VGND VGND VPWR VPWR _12776_/X sky130_fd_sc_hd__o22a_1
X_15564_ _15566_/CLK _15564_/D VGND VGND VPWR VPWR _15564_/Q sky130_fd_sc_hd__dfxtp_2
X_14515_ _11632_/X _14515_/D VGND VGND VPWR VPWR _14515_/Q sky130_fd_sc_hd__dfxtp_1
X_11727_ _11731_/A VGND VGND VPWR VPWR _11727_/X sky130_fd_sc_hd__clkbuf_1
X_15495_ _15591_/CLK _15495_/D VGND VGND VPWR VPWR wdata[21] sky130_fd_sc_hd__dfxtp_2
X_14446_ _11871_/X _14446_/D VGND VGND VPWR VPWR _14446_/Q sky130_fd_sc_hd__dfxtp_1
X_11658_ _11658_/A VGND VGND VPWR VPWR _11658_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10609_ _14771_/Q _10607_/X _10367_/X _10608_/X VGND VGND VPWR VPWR _14771_/D sky130_fd_sc_hd__a22o_1
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ _14385_/CLK instruction[6] VGND VGND VPWR VPWR _14377_/Q sky130_fd_sc_hd__dfxtp_2
X_11589_ _11589_/A VGND VGND VPWR VPWR _11651_/A sky130_fd_sc_hd__buf_2
X_13328_ _13331_/X _13329_/X _13393_/S VGND VGND VPWR VPWR _13328_/X sky130_fd_sc_hd__mux2_2
XFILLER_115_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13259_ _12737_/A _12758_/A _13418_/S VGND VGND VPWR VPWR _13259_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07820_ _07820_/A _07820_/B _07820_/C VGND VGND VPWR VPWR _15451_/D sky130_fd_sc_hd__and3_1
XFILLER_97_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07751_ _07748_/X _07750_/X _07748_/X _07750_/X VGND VGND VPWR VPWR _07895_/B sky130_fd_sc_hd__a2bb2o_1
X_07682_ _07689_/A VGND VGND VPWR VPWR _07682_/X sky130_fd_sc_hd__buf_1
XFILLER_65_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09421_ _15072_/Q _09410_/X _09164_/X _09413_/X VGND VGND VPWR VPWR _15072_/D sky130_fd_sc_hd__a22o_1
X_09352_ _15092_/Q _09345_/X _09220_/X _09347_/X VGND VGND VPWR VPWR _15092_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08303_ _15342_/Q _08291_/X _08042_/X _08292_/X VGND VGND VPWR VPWR _15342_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09283_ _09289_/A VGND VGND VPWR VPWR _09283_/X sky130_fd_sc_hd__buf_1
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08234_ _08238_/A VGND VGND VPWR VPWR _08234_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08165_ _08174_/A VGND VGND VPWR VPWR _08165_/X sky130_fd_sc_hd__buf_1
XFILLER_107_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07116_ _07835_/A VGND VGND VPWR VPWR _07820_/A sky130_fd_sc_hd__buf_1
XFILLER_118_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08096_ _15396_/Q _07927_/A _08095_/X _07932_/A VGND VGND VPWR VPWR _15396_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08998_ _08998_/A VGND VGND VPWR VPWR _08998_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07949_ _07981_/A VGND VGND VPWR VPWR _07949_/X sky130_fd_sc_hd__buf_1
XFILLER_29_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10960_ _14688_/Q _10951_/X _10677_/X _10954_/X VGND VGND VPWR VPWR _14688_/D sky130_fd_sc_hd__a22o_1
XFILLER_44_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09619_ _09634_/A VGND VGND VPWR VPWR _09630_/A sky130_fd_sc_hd__buf_1
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10891_ _14708_/Q _10884_/X _10746_/X _10886_/X VGND VGND VPWR VPWR _14708_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12630_ _12946_/A _12091_/X _12360_/A VGND VGND VPWR VPWR _12632_/A sky130_fd_sc_hd__o21ai_1
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _12561_/A _12561_/B VGND VGND VPWR VPWR _12561_/Y sky130_fd_sc_hd__nor2_1
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11512_ _11517_/A VGND VGND VPWR VPWR _11512_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14300_ _15469_/CLK _15467_/Q VGND VGND VPWR VPWR _14300_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15280_ _08616_/X _15280_/D VGND VGND VPWR VPWR _15280_/Q sky130_fd_sc_hd__dfxtp_1
X_12492_ _12492_/A VGND VGND VPWR VPWR _12492_/X sky130_fd_sc_hd__clkbuf_4
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ _14227_/X _14228_/X _14229_/X _14230_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14231_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11443_ _11443_/A VGND VGND VPWR VPWR _11443_/X sky130_fd_sc_hd__buf_1
XFILLER_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14162_ _15215_/Q _14543_/Q _14991_/Q _15407_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14162_/X sky130_fd_sc_hd__mux4_2
XFILLER_152_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11374_ _11384_/A VGND VGND VPWR VPWR _11374_/X sky130_fd_sc_hd__buf_1
XFILLER_124_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13113_ _15659_/Q data_address[24] _15667_/Q VGND VGND VPWR VPWR _13113_/X sky130_fd_sc_hd__mux2_1
X_10325_ _14845_/Q _10313_/X _10324_/X _10317_/X VGND VGND VPWR VPWR _14845_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14093_ _14678_/Q _15254_/Q _14742_/Q _14710_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14093_/X sky130_fd_sc_hd__mux4_2
XFILLER_79_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13044_ wdata[17] rdata[17] ren VGND VGND VPWR VPWR _14321_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10256_ _10256_/A VGND VGND VPWR VPWR _10280_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10187_ _14882_/Q _10183_/X _09928_/X _10186_/X VGND VGND VPWR VPWR _14882_/D sky130_fd_sc_hd__a22o_1
XFILLER_121_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14995_ _09755_/X _14995_/D VGND VGND VPWR VPWR _14995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13946_ _13942_/X _13943_/X _13944_/X _13945_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13946_/X sky130_fd_sc_hd__mux4_2
XFILLER_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13877_ _14636_/Q _14604_/Q _14572_/Q _15372_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13877_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15616_ _15647_/CLK _15616_/D VGND VGND VPWR VPWR pc[11] sky130_fd_sc_hd__dfxtp_2
X_12828_ _15535_/Q VGND VGND VPWR VPWR _12828_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15547_ _15566_/CLK _15547_/D VGND VGND VPWR VPWR _15547_/Q sky130_fd_sc_hd__dfxtp_1
X_12759_ _13267_/X _12698_/X _13262_/X _12701_/X _12758_/X VGND VGND VPWR VPWR _12759_/X
+ sky130_fd_sc_hd__o221a_1
X_15478_ _15509_/CLK _15478_/D VGND VGND VPWR VPWR wdata[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_147_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14429_ _11932_/X _14429_/D VGND VGND VPWR VPWR _14429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09970_ _14938_/Q _09957_/X _09969_/X _09959_/X VGND VGND VPWR VPWR _14938_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08921_ _08921_/A VGND VGND VPWR VPWR _08936_/A sky130_fd_sc_hd__buf_1
XFILLER_130_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08852_ _09224_/A VGND VGND VPWR VPWR _08852_/X sky130_fd_sc_hd__buf_1
XFILLER_85_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07803_ _07803_/A VGND VGND VPWR VPWR _07805_/A sky130_fd_sc_hd__inv_2
XFILLER_84_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08783_ _09153_/A VGND VGND VPWR VPWR _08783_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_49_clk _14315_/CLK VGND VGND VPWR VPWR _15669_/CLK sky130_fd_sc_hd__clkbuf_16
X_07734_ _07723_/X _07725_/X _07720_/Y _13141_/X _07679_/A VGND VGND VPWR VPWR _07734_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07665_ _07663_/X _07664_/X _07663_/X _13124_/X VGND VGND VPWR VPWR _07798_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09404_ _15076_/Q _09298_/A _09287_/X _09301_/A VGND VGND VPWR VPWR _15076_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07596_ _07596_/A VGND VGND VPWR VPWR _07599_/A sky130_fd_sc_hd__buf_1
XFILLER_80_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09335_ _09335_/A VGND VGND VPWR VPWR _09335_/X sky130_fd_sc_hd__buf_1
X_09266_ _09266_/A VGND VGND VPWR VPWR _09266_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08217_ _14302_/Q VGND VGND VPWR VPWR _09923_/B sky130_fd_sc_hd__inv_2
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09197_ _09197_/A VGND VGND VPWR VPWR _09197_/X sky130_fd_sc_hd__buf_1
XFILLER_153_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08148_ _08148_/A VGND VGND VPWR VPWR _08148_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08079_ _08079_/A VGND VGND VPWR VPWR _08079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10110_ _14904_/Q _10106_/X _09977_/X _10107_/X VGND VGND VPWR VPWR _14904_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11090_ _11098_/A VGND VGND VPWR VPWR _11090_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10041_ _10041_/A VGND VGND VPWR VPWR _10041_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13800_ _14964_/Q _15060_/Q _15028_/Q _15092_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13800_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11992_ _11992_/A VGND VGND VPWR VPWR _11992_/X sky130_fd_sc_hd__clkbuf_1
X_14780_ _10574_/X _14780_/D VGND VGND VPWR VPWR _14780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10943_ _10956_/A VGND VGND VPWR VPWR _10948_/A sky130_fd_sc_hd__buf_1
X_13731_ _13727_/X _13728_/X _13729_/X _13730_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13731_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10874_ _10874_/A VGND VGND VPWR VPWR _10874_/X sky130_fd_sc_hd__buf_1
X_13662_ _15233_/Q _14561_/Q _15009_/Q _15425_/Q _13740_/S0 _07541_/A VGND VGND VPWR
+ VPWR _13662_/X sky130_fd_sc_hd__mux4_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15401_ _08067_/X _15401_/D VGND VGND VPWR VPWR _15401_/Q sky130_fd_sc_hd__dfxtp_1
X_12613_ _12611_/X _12097_/A _12612_/Y VGND VGND VPWR VPWR _12613_/X sky130_fd_sc_hd__o21a_1
X_13593_ _13592_/X _07310_/Y _13649_/S VGND VGND VPWR VPWR _13593_/X sky130_fd_sc_hd__mux2_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12544_ _15473_/Q VGND VGND VPWR VPWR _12545_/C sky130_fd_sc_hd__inv_2
X_15332_ _08334_/X _15332_/D VGND VGND VPWR VPWR _15332_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15263_ _08676_/X _15263_/D VGND VGND VPWR VPWR _15263_/Q sky130_fd_sc_hd__dfxtp_1
X_12475_ _12727_/A VGND VGND VPWR VPWR _12475_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11426_ _14563_/Q _11319_/A _11201_/X _11322_/A VGND VGND VPWR VPWR _14563_/D sky130_fd_sc_hd__a22o_1
X_14214_ _15178_/Q _15146_/Q _14762_/Q _14794_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14214_/X sky130_fd_sc_hd__mux4_1
X_15194_ _08959_/X _15194_/D VGND VGND VPWR VPWR _15194_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_6 data_address[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14145_ _15121_/Q _15345_/Q _15313_/Q _15281_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14145_/X sky130_fd_sc_hd__mux4_2
X_11357_ _11368_/A VGND VGND VPWR VPWR _11362_/A sky130_fd_sc_hd__buf_2
X_10308_ _10308_/A VGND VGND VPWR VPWR _10308_/X sky130_fd_sc_hd__buf_1
X_14076_ _14072_/X _14073_/X _14074_/X _14075_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14076_/X sky130_fd_sc_hd__mux4_2
XFILLER_113_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11288_ _11290_/A VGND VGND VPWR VPWR _11288_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13027_ wdata[0] rdata[0] _13058_/S VGND VGND VPWR VPWR _14304_/D sky130_fd_sc_hd__mux2_1
X_10239_ _14867_/Q _10237_/X _09999_/X _10238_/X VGND VGND VPWR VPWR _14867_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14978_ _09809_/X _14978_/D VGND VGND VPWR VPWR _14978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13929_ _14823_/Q _14855_/Q _14887_/Q _14919_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13929_/X sky130_fd_sc_hd__mux4_1
X_07450_ _07451_/A _13442_/X VGND VGND VPWR VPWR _15556_/D sky130_fd_sc_hd__and2_1
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07381_ _13156_/X _07363_/X _07509_/B _07319_/A _07380_/X VGND VGND VPWR VPWR _07385_/B
+ sky130_fd_sc_hd__o221a_2
X_09120_ _09120_/A VGND VGND VPWR VPWR _09125_/A sky130_fd_sc_hd__buf_1
XFILLER_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09051_ _09051_/A VGND VGND VPWR VPWR _09051_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08002_ _08032_/A VGND VGND VPWR VPWR _08002_/X sky130_fd_sc_hd__buf_1
XFILLER_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09953_ _09961_/A VGND VGND VPWR VPWR _09953_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08904_ _08904_/A VGND VGND VPWR VPWR _08904_/X sky130_fd_sc_hd__buf_1
XFILLER_131_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09884_ _14958_/Q _09877_/X _09637_/X _09878_/X VGND VGND VPWR VPWR _14958_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08835_ _15223_/Q _08825_/X _08834_/X _08827_/X VGND VGND VPWR VPWR _15223_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08766_ _08770_/A VGND VGND VPWR VPWR _08766_/X sky130_fd_sc_hd__clkbuf_1
X_07717_ _07715_/X _13139_/X _07710_/X VGND VGND VPWR VPWR _07868_/A sky130_fd_sc_hd__a21bo_1
X_08697_ _08701_/A VGND VGND VPWR VPWR _08697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07648_ _07687_/A VGND VGND VPWR VPWR _07701_/A sky130_fd_sc_hd__buf_1
XFILLER_81_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07579_ _07581_/A _13082_/X VGND VGND VPWR VPWR _15497_/D sky130_fd_sc_hd__and2_1
X_09318_ _09318_/A VGND VGND VPWR VPWR _09318_/X sky130_fd_sc_hd__clkbuf_1
X_10590_ _10610_/A VGND VGND VPWR VPWR _10595_/A sky130_fd_sc_hd__buf_2
X_09249_ _09274_/A VGND VGND VPWR VPWR _09249_/X sky130_fd_sc_hd__buf_1
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12260_ _15533_/Q VGND VGND VPWR VPWR _12854_/A sky130_fd_sc_hd__buf_1
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11211_ _14626_/Q _11207_/X _11065_/X _11210_/X VGND VGND VPWR VPWR _14626_/D sky130_fd_sc_hd__a22o_1
X_12191_ _12750_/A VGND VGND VPWR VPWR _12191_/Y sky130_fd_sc_hd__inv_2
X_11142_ _11168_/A VGND VGND VPWR VPWR _11151_/A sky130_fd_sc_hd__buf_1
XFILLER_150_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11073_ _11089_/A VGND VGND VPWR VPWR _11086_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14901_ _10121_/X _14901_/D VGND VGND VPWR VPWR _14901_/Q sky130_fd_sc_hd__dfxtp_1
X_10024_ _10050_/A VGND VGND VPWR VPWR _10024_/X sky130_fd_sc_hd__buf_1
XFILLER_49_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14832_ _10377_/X _14832_/D VGND VGND VPWR VPWR _14832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14763_ _10634_/X _14763_/D VGND VGND VPWR VPWR _14763_/Q sky130_fd_sc_hd__dfxtp_1
X_11975_ _11981_/A VGND VGND VPWR VPWR _11975_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13714_ _15196_/Q _15164_/Q _14780_/Q _14812_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13714_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10926_ _14698_/Q _10924_/X _10799_/X _10925_/X VGND VGND VPWR VPWR _14698_/D sky130_fd_sc_hd__a22o_1
X_14694_ _10939_/X _14694_/D VGND VGND VPWR VPWR _14694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10857_ _14719_/Q _10853_/X _10684_/X _10856_/X VGND VGND VPWR VPWR _14719_/D sky130_fd_sc_hd__a22o_1
X_13645_ _13644_/X _07382_/Y _13649_/S VGND VGND VPWR VPWR _13645_/X sky130_fd_sc_hd__mux2_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _14106_/X _14111_/X _13648_/S VGND VGND VPWR VPWR _13576_/X sky130_fd_sc_hd__mux2_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ _11533_/A VGND VGND VPWR VPWR _10788_/X sky130_fd_sc_hd__buf_1
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15315_ _08444_/X _15315_/D VGND VGND VPWR VPWR _15315_/Q sky130_fd_sc_hd__dfxtp_1
X_12527_ _12962_/A _12522_/X _12502_/X VGND VGND VPWR VPWR _12527_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15246_ _08738_/X _15246_/D VGND VGND VPWR VPWR _15246_/Q sky130_fd_sc_hd__dfxtp_1
X_12458_ _12819_/A _13363_/X VGND VGND VPWR VPWR _12459_/B sky130_fd_sc_hd__or2_1
X_11409_ _11413_/A VGND VGND VPWR VPWR _11409_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12389_ _12452_/A VGND VGND VPWR VPWR _12389_/X sky130_fd_sc_hd__buf_1
X_15177_ _09019_/X _15177_/D VGND VGND VPWR VPWR _15177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14128_ _14515_/Q _14483_/Q _14451_/Q _14419_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14128_/X sky130_fd_sc_hd__mux4_2
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14059_ _14842_/Q _14874_/Q _14906_/Q _14938_/Q _14395_/Q _14060_/S1 VGND VGND VPWR
+ VPWR _14059_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08620_ _08622_/A VGND VGND VPWR VPWR _08620_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08551_ _08563_/A VGND VGND VPWR VPWR _08552_/A sky130_fd_sc_hd__buf_1
XFILLER_82_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07502_ _07511_/A VGND VGND VPWR VPWR _07506_/A sky130_fd_sc_hd__buf_1
X_08482_ _08520_/A VGND VGND VPWR VPWR _08482_/X sky130_fd_sc_hd__buf_1
XFILLER_63_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07433_ _07473_/A VGND VGND VPWR VPWR _07460_/A sky130_fd_sc_hd__buf_1
XFILLER_23_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07364_ _14381_/Q VGND VGND VPWR VPWR _07508_/B sky130_fd_sc_hd__inv_2
XFILLER_149_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09103_ _09105_/A VGND VGND VPWR VPWR _09103_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07295_ _14374_/Q _14373_/Q _14372_/Q _14371_/Q VGND VGND VPWR VPWR _07559_/B sky130_fd_sc_hd__or4bb_4
XFILLER_108_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09034_ _09038_/A VGND VGND VPWR VPWR _09034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09936_ _09952_/A VGND VGND VPWR VPWR _09949_/A sky130_fd_sc_hd__buf_1
X_09867_ _09867_/A VGND VGND VPWR VPWR _09867_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08818_ _15227_/Q _08812_/X _08817_/X _08814_/X VGND VGND VPWR VPWR _15227_/D sky130_fd_sc_hd__a22o_1
X_09798_ _09798_/A VGND VGND VPWR VPWR _09798_/X sky130_fd_sc_hd__buf_1
XANTENNA_204 _13570_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08749_ _15244_/Q _08742_/X _08492_/X _08744_/X VGND VGND VPWR VPWR _15244_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_215 _13462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_226 _08588_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_237 _11216_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11760_ _11762_/A VGND VGND VPWR VPWR _11760_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_248 _11900_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_259 _14314_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10711_ _10721_/A VGND VGND VPWR VPWR _10711_/X sky130_fd_sc_hd__clkbuf_1
X_11691_ _11691_/A VGND VGND VPWR VPWR _11691_/X sky130_fd_sc_hd__buf_1
XFILLER_14_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13430_ _13429_/X _13090_/X _14336_/Q VGND VGND VPWR VPWR _13430_/X sky130_fd_sc_hd__mux2_1
X_10642_ _14761_/Q _10637_/X _10411_/X _10638_/X VGND VGND VPWR VPWR _14761_/D sky130_fd_sc_hd__a22o_1
XFILLER_10_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13361_ _13368_/X _13362_/X _13393_/S VGND VGND VPWR VPWR _13361_/X sky130_fd_sc_hd__mux2_2
X_10573_ _14781_/Q _10564_/X _10324_/X _10567_/X VGND VGND VPWR VPWR _14781_/D sky130_fd_sc_hd__a22o_1
X_15100_ _09325_/X _15100_/D VGND VGND VPWR VPWR _15100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12312_ _12663_/A VGND VGND VPWR VPWR _12745_/A sky130_fd_sc_hd__buf_2
X_13292_ _13293_/X _12521_/B _13393_/S VGND VGND VPWR VPWR _13292_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12243_ _15567_/Q VGND VGND VPWR VPWR _12243_/X sky130_fd_sc_hd__clkbuf_2
X_15031_ _09587_/X _15031_/D VGND VGND VPWR VPWR _15031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12174_ _12172_/X _12082_/X _12726_/A _12084_/X VGND VGND VPWR VPWR _12271_/B sky130_fd_sc_hd__o22a_1
XFILLER_122_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11125_ _11125_/A VGND VGND VPWR VPWR _11125_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11056_ _11101_/A VGND VGND VPWR VPWR _11089_/A sky130_fd_sc_hd__clkbuf_2
X_10007_ _10015_/A VGND VGND VPWR VPWR _10007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14815_ _10450_/X _14815_/D VGND VGND VPWR VPWR _14815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14746_ _10711_/X _14746_/D VGND VGND VPWR VPWR _14746_/Q sky130_fd_sc_hd__dfxtp_1
X_11958_ _11977_/A VGND VGND VPWR VPWR _11958_/X sky130_fd_sc_hd__buf_1
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10909_ _10909_/A VGND VGND VPWR VPWR _10909_/X sky130_fd_sc_hd__clkbuf_1
X_14677_ _11001_/X _14677_/D VGND VGND VPWR VPWR _14677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11889_ _11889_/A VGND VGND VPWR VPWR _11889_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater40 _14238_/S1 VGND VGND VPWR VPWR _07379_/A sky130_fd_sc_hd__clkbuf_16
X_13628_ _14236_/X _14241_/X _13648_/S VGND VGND VPWR VPWR _13628_/X sky130_fd_sc_hd__mux2_2
Xrepeater51 _14395_/Q VGND VGND VPWR VPWR _14060_/S0 sky130_fd_sc_hd__clkbuf_16
XFILLER_32_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13559_ _13558_/X _13082_/X _14337_/Q VGND VGND VPWR VPWR _13559_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15229_ _08808_/X _15229_/D VGND VGND VPWR VPWR _15229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07982_ _14326_/Q VGND VGND VPWR VPWR _07983_/A sky130_fd_sc_hd__buf_1
X_09721_ _15006_/Q _09715_/X _09553_/X _09718_/X VGND VGND VPWR VPWR _15006_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09652_ _09860_/A VGND VGND VPWR VPWR _09733_/A sky130_fd_sc_hd__buf_1
XFILLER_67_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08603_ _08603_/A VGND VGND VPWR VPWR _08603_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09583_ _10722_/A VGND VGND VPWR VPWR _10344_/A sky130_fd_sc_hd__buf_1
XFILLER_103_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08534_ _10823_/A VGND VGND VPWR VPWR _09284_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08465_ _10765_/A VGND VGND VPWR VPWR _09236_/A sky130_fd_sc_hd__clkbuf_2
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07416_ _07416_/A VGND VGND VPWR VPWR _07419_/A sky130_fd_sc_hd__buf_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08396_ _09188_/A VGND VGND VPWR VPWR _08396_/X sky130_fd_sc_hd__buf_1
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07347_ _07495_/B _07339_/X _07497_/B _07341_/X VGND VGND VPWR VPWR _07349_/B sky130_fd_sc_hd__o22a_1
XFILLER_109_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07278_ _07278_/A _07278_/B VGND VGND VPWR VPWR _15616_/D sky130_fd_sc_hd__nor2_1
XFILLER_124_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09017_ _09026_/A VGND VGND VPWR VPWR _09017_/X sky130_fd_sc_hd__buf_1
XFILLER_88_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09919_ _09933_/A VGND VGND VPWR VPWR _09919_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12930_ _12213_/Y _12867_/B _12957_/C _12928_/X _12929_/X VGND VGND VPWR VPWR _12930_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_46_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12861_ _12861_/A VGND VGND VPWR VPWR _12861_/X sky130_fd_sc_hd__buf_1
XFILLER_73_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14600_ _11299_/X _14600_/D VGND VGND VPWR VPWR _14600_/Q sky130_fd_sc_hd__dfxtp_1
X_11812_ _11874_/A VGND VGND VPWR VPWR _11834_/A sky130_fd_sc_hd__buf_2
X_15580_ _15592_/CLK _15580_/D VGND VGND VPWR VPWR _15580_/Q sky130_fd_sc_hd__dfxtp_1
X_12792_ _12775_/X _12788_/X _12715_/X VGND VGND VPWR VPWR _12792_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14531_ _11569_/X _14531_/D VGND VGND VPWR VPWR _14531_/Q sky130_fd_sc_hd__dfxtp_1
X_11743_ _11752_/A VGND VGND VPWR VPWR _11743_/X sky130_fd_sc_hd__buf_1
XFILLER_42_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14462_ _11818_/X _14462_/D VGND VGND VPWR VPWR _14462_/Q sky130_fd_sc_hd__dfxtp_1
X_11674_ _11674_/A VGND VGND VPWR VPWR _11674_/X sky130_fd_sc_hd__buf_1
XFILLER_41_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13413_ _12762_/X _12758_/A _13418_/S VGND VGND VPWR VPWR _13413_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10625_ _10625_/A VGND VGND VPWR VPWR _10625_/X sky130_fd_sc_hd__clkbuf_1
X_14393_ _14393_/CLK instruction[30] VGND VGND VPWR VPWR _14393_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13344_ _13347_/X _13345_/X _13393_/S VGND VGND VPWR VPWR _13344_/X sky130_fd_sc_hd__mux2_1
X_10556_ _10578_/A VGND VGND VPWR VPWR _10561_/A sky130_fd_sc_hd__buf_1
XFILLER_143_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13275_ _13276_/X _13305_/X _15563_/Q VGND VGND VPWR VPWR _13275_/X sky130_fd_sc_hd__mux2_1
X_10487_ _14806_/Q _10484_/X _10354_/X _10486_/X VGND VGND VPWR VPWR _14806_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15014_ _09680_/X _15014_/D VGND VGND VPWR VPWR _15014_/Q sky130_fd_sc_hd__dfxtp_1
X_12226_ _12223_/A _12225_/X _12223_/A _12225_/X VGND VGND VPWR VPWR _12892_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12157_ _12157_/A VGND VGND VPWR VPWR _12157_/X sky130_fd_sc_hd__buf_1
XFILLER_123_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11108_ _11475_/A VGND VGND VPWR VPWR _11108_/X sky130_fd_sc_hd__buf_1
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12088_ _12588_/A _12087_/B _12087_/Y VGND VGND VPWR VPWR _12585_/A sky130_fd_sc_hd__a21oi_4
XFILLER_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11039_ _14666_/Q _11037_/X _10799_/X _11038_/X VGND VGND VPWR VPWR _14666_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14729_ _10802_/X _14729_/D VGND VGND VPWR VPWR _14729_/Q sky130_fd_sc_hd__dfxtp_1
X_08250_ _15357_/Q _08241_/X _07963_/X _08244_/X VGND VGND VPWR VPWR _15357_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07201_ _07259_/B _07173_/B _07200_/X _07197_/Y VGND VGND VPWR VPWR _15659_/D sky130_fd_sc_hd__a211oi_4
XFILLER_20_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08181_ _08189_/A VGND VGND VPWR VPWR _08181_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07132_ _13112_/X VGND VGND VPWR VPWR _07260_/B sky130_fd_sc_hd__inv_2
XFILLER_118_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07965_ _07971_/A VGND VGND VPWR VPWR _07965_/X sky130_fd_sc_hd__clkbuf_1
X_09704_ _09716_/A VGND VGND VPWR VPWR _09705_/A sky130_fd_sc_hd__buf_1
XFILLER_114_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07896_ _07748_/X _07750_/X _07895_/X VGND VGND VPWR VPWR _07897_/B sky130_fd_sc_hd__o21ai_1
XFILLER_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09635_ _09647_/A VGND VGND VPWR VPWR _09635_/X sky130_fd_sc_hd__buf_1
XFILLER_43_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09566_ _15036_/Q _09562_/X _09564_/X _09565_/X VGND VGND VPWR VPWR _15036_/D sky130_fd_sc_hd__a22o_1
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ _09271_/A VGND VGND VPWR VPWR _08517_/X sky130_fd_sc_hd__buf_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09497_ _09506_/A VGND VGND VPWR VPWR _09497_/X sky130_fd_sc_hd__buf_1
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08448_ _09224_/A VGND VGND VPWR VPWR _08448_/X sky130_fd_sc_hd__buf_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08379_ _08379_/A VGND VGND VPWR VPWR _08416_/A sky130_fd_sc_hd__buf_1
XFILLER_7_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10410_ _10410_/A VGND VGND VPWR VPWR _10410_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11390_ _11392_/A VGND VGND VPWR VPWR _11390_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10341_ _10341_/A VGND VGND VPWR VPWR _10341_/X sky130_fd_sc_hd__buf_1
XFILLER_136_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13060_ _12894_/Y _15562_/Q _13076_/S VGND VGND VPWR VPWR _13060_/X sky130_fd_sc_hd__mux2_1
X_10272_ _10492_/A VGND VGND VPWR VPWR _10346_/A sky130_fd_sc_hd__buf_1
XFILLER_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12011_ _14405_/Q _12005_/X _08091_/A _12006_/X VGND VGND VPWR VPWR _14405_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13962_ _15203_/Q _14531_/Q _14979_/Q _15395_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13962_/X sky130_fd_sc_hd__mux4_2
XFILLER_93_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12913_ _12913_/A _12913_/B VGND VGND VPWR VPWR _12913_/X sky130_fd_sc_hd__or2_1
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13893_ _14666_/Q _15242_/Q _14730_/Q _14698_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13893_/X sky130_fd_sc_hd__mux4_2
X_15632_ _15663_/CLK _15632_/D VGND VGND VPWR VPWR pc[27] sky130_fd_sc_hd__dfxtp_4
X_12844_ _12847_/A _12847_/B _12328_/X VGND VGND VPWR VPWR _12844_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15563_ _15566_/CLK _15563_/D VGND VGND VPWR VPWR _15563_/Q sky130_fd_sc_hd__dfxtp_4
X_12775_ _12775_/A VGND VGND VPWR VPWR _12775_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14514_ _11636_/X _14514_/D VGND VGND VPWR VPWR _14514_/Q sky130_fd_sc_hd__dfxtp_1
X_11726_ _11746_/A VGND VGND VPWR VPWR _11731_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15494_ _15579_/CLK _15494_/D VGND VGND VPWR VPWR wdata[20] sky130_fd_sc_hd__dfxtp_4
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14445_ _11873_/X _14445_/D VGND VGND VPWR VPWR _14445_/Q sky130_fd_sc_hd__dfxtp_1
X_11657_ _14508_/Q _11652_/X _11533_/X _11654_/X VGND VGND VPWR VPWR _14508_/D sky130_fd_sc_hd__a22o_1
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10608_ _10617_/A VGND VGND VPWR VPWR _10608_/X sky130_fd_sc_hd__buf_1
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _14385_/CLK instruction[5] VGND VGND VPWR VPWR _14376_/Q sky130_fd_sc_hd__dfxtp_2
X_11588_ _11598_/A VGND VGND VPWR VPWR _11588_/X sky130_fd_sc_hd__clkbuf_1
X_13327_ _13326_/X _13328_/X _15565_/Q VGND VGND VPWR VPWR _13327_/X sky130_fd_sc_hd__mux2_1
X_10539_ _14790_/Q _10535_/X _10423_/X _10536_/X VGND VGND VPWR VPWR _14790_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13258_ _13259_/X _13271_/X _13415_/S VGND VGND VPWR VPWR _13258_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12209_ _12209_/A _12209_/B _12746_/A VGND VGND VPWR VPWR _12209_/X sky130_fd_sc_hd__or3b_1
XFILLER_151_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13189_ _13188_/X _13230_/X _13393_/S VGND VGND VPWR VPWR _13189_/X sky130_fd_sc_hd__mux2_1
X_07750_ _07766_/B VGND VGND VPWR VPWR _07750_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07681_ _07706_/A _13135_/X VGND VGND VPWR VPWR _07681_/X sky130_fd_sc_hd__or2_1
XFILLER_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09420_ _09422_/A VGND VGND VPWR VPWR _09420_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09351_ _09351_/A VGND VGND VPWR VPWR _09351_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08302_ _08304_/A VGND VGND VPWR VPWR _08302_/X sky130_fd_sc_hd__clkbuf_1
X_09282_ _09307_/A VGND VGND VPWR VPWR _09289_/A sky130_fd_sc_hd__buf_1
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08233_ _08255_/A VGND VGND VPWR VPWR _08238_/A sky130_fd_sc_hd__buf_1
XFILLER_119_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08164_ _08173_/A VGND VGND VPWR VPWR _08164_/X sky130_fd_sc_hd__buf_1
XFILLER_119_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07115_ _07795_/A VGND VGND VPWR VPWR _07835_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_146_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08095_ _08095_/A VGND VGND VPWR VPWR _08095_/X sky130_fd_sc_hd__buf_1
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08997_ _15183_/Q _08993_/X _08869_/X _08994_/X VGND VGND VPWR VPWR _15183_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07948_ _08045_/A VGND VGND VPWR VPWR _07981_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07879_ _07723_/X _07725_/X _07878_/Y VGND VGND VPWR VPWR _07880_/A sky130_fd_sc_hd__o21ai_1
XFILLER_83_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09618_ _15026_/Q _09610_/X _09617_/X _09613_/X VGND VGND VPWR VPWR _15026_/D sky130_fd_sc_hd__a22o_1
X_10890_ _10890_/A VGND VGND VPWR VPWR _10890_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09549_ _09580_/A VGND VGND VPWR VPWR _09549_/X sky130_fd_sc_hd__buf_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12560_ _12546_/X _12559_/Y _12553_/X VGND VGND VPWR VPWR wstrobe[2] sky130_fd_sc_hd__o21a_4
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11511_ _14545_/Q _11501_/X _11510_/X _11503_/X VGND VGND VPWR VPWR _14545_/D sky130_fd_sc_hd__a22o_1
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12491_/A VGND VGND VPWR VPWR _12492_/A sky130_fd_sc_hd__buf_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14230_ _14953_/Q _15049_/Q _15017_/Q _15081_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14230_/X sky130_fd_sc_hd__mux4_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11442_ _11454_/A VGND VGND VPWR VPWR _11442_/X sky130_fd_sc_hd__buf_1
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14161_ _14157_/X _14158_/X _14159_/X _14160_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14161_/X sky130_fd_sc_hd__mux4_1
X_11373_ _11373_/A VGND VGND VPWR VPWR _11373_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13112_ _15658_/Q data_address[23] _15667_/Q VGND VGND VPWR VPWR _13112_/X sky130_fd_sc_hd__mux2_1
X_10324_ _10324_/A VGND VGND VPWR VPWR _10324_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14092_ _15222_/Q _14550_/Q _14998_/Q _15414_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14092_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13043_ wdata[16] rdata[16] ren VGND VGND VPWR VPWR _14320_/D sky130_fd_sc_hd__mux2_1
X_10255_ _10255_/A VGND VGND VPWR VPWR _10255_/X sky130_fd_sc_hd__buf_1
XFILLER_152_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10186_ _10186_/A VGND VGND VPWR VPWR _10186_/X sky130_fd_sc_hd__buf_1
X_14994_ _09759_/X _14994_/D VGND VGND VPWR VPWR _14994_/Q sky130_fd_sc_hd__dfxtp_1
X_13945_ _15109_/Q _15333_/Q _15301_/Q _15269_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13945_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13876_ _13872_/X _13873_/X _13874_/X _13875_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13876_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15615_ _15647_/CLK _15615_/D VGND VGND VPWR VPWR pc[10] sky130_fd_sc_hd__dfxtp_4
XFILLER_61_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12827_ _12820_/X _12825_/X _12789_/X _13300_/X _12826_/X VGND VGND VPWR VPWR _12827_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_50_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15546_ _15566_/CLK _15546_/D VGND VGND VPWR VPWR _15546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12758_ _12758_/A _12758_/B _12758_/C VGND VGND VPWR VPWR _12758_/X sky130_fd_sc_hd__or3_2
XFILLER_61_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11709_ _14494_/Q _11702_/X _11455_/X _11705_/X VGND VGND VPWR VPWR _14494_/D sky130_fd_sc_hd__a22o_1
X_15477_ _15521_/CLK _15477_/D VGND VGND VPWR VPWR wdata[3] sky130_fd_sc_hd__dfxtp_2
X_12689_ _12689_/A _12689_/B VGND VGND VPWR VPWR _12690_/B sky130_fd_sc_hd__nand2_2
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14428_ _11935_/X _14428_/D VGND VGND VPWR VPWR _14428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14359_ _15654_/CLK pc[20] VGND VGND VPWR VPWR _14359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08920_ _15203_/Q _08782_/A _08919_/X _08786_/A VGND VGND VPWR VPWR _15203_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08851_ _08864_/A VGND VGND VPWR VPWR _08851_/X sky130_fd_sc_hd__buf_1
XFILLER_112_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07802_ _07785_/Y _07666_/Y _07796_/X _07798_/X VGND VGND VPWR VPWR _15455_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08782_ _08782_/A VGND VGND VPWR VPWR _08782_/X sky130_fd_sc_hd__buf_1
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07733_ _07733_/A VGND VGND VPWR VPWR _07733_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07664_ _13124_/X VGND VGND VPWR VPWR _07664_/X sky130_fd_sc_hd__buf_1
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09403_ _09407_/A VGND VGND VPWR VPWR _09403_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07595_ _07595_/A _13071_/X VGND VGND VPWR VPWR _15486_/D sky130_fd_sc_hd__and2_1
XFILLER_53_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09334_ _09340_/A VGND VGND VPWR VPWR _09334_/X sky130_fd_sc_hd__clkbuf_1
X_09265_ _15114_/Q _09262_/X _09263_/X _09264_/X VGND VGND VPWR VPWR _15114_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08216_ _08216_/A VGND VGND VPWR VPWR _08216_/X sky130_fd_sc_hd__clkbuf_1
X_09196_ _09196_/A VGND VGND VPWR VPWR _09196_/X sky130_fd_sc_hd__buf_1
XFILLER_5_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08147_ _15384_/Q _08143_/X _07988_/X _08144_/X VGND VGND VPWR VPWR _15384_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08078_ _14308_/Q VGND VGND VPWR VPWR _08079_/A sky130_fd_sc_hd__buf_1
XFILLER_1_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10040_ _14922_/Q _10037_/X _10038_/X _10039_/X VGND VGND VPWR VPWR _14922_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11991_ _14412_/Q _11986_/X _08054_/A _11988_/X VGND VGND VPWR VPWR _14412_/D sky130_fd_sc_hd__a22o_1
XFILLER_72_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13730_ _14971_/Q _15067_/Q _15035_/Q _15099_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13730_/X sky130_fd_sc_hd__mux4_1
X_10942_ _14693_/Q _10936_/X _10824_/X _10937_/X VGND VGND VPWR VPWR _14693_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13661_ _13657_/X _13658_/X _13659_/X _13660_/X _07533_/A _14402_/Q VGND VGND VPWR
+ VPWR _13661_/X sky130_fd_sc_hd__mux4_1
X_10873_ _10879_/A VGND VGND VPWR VPWR _10873_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15400_ _08072_/X _15400_/D VGND VGND VPWR VPWR _15400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12612_ _12625_/A _12625_/B VGND VGND VPWR VPWR _12612_/Y sky130_fd_sc_hd__nand2_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13592_ _14146_/X _14151_/X _13648_/S VGND VGND VPWR VPWR _13592_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15331_ _08337_/X _15331_/D VGND VGND VPWR VPWR _15331_/Q sky130_fd_sc_hd__dfxtp_1
X_12543_ _15472_/Q VGND VGND VPWR VPWR _12551_/A sky130_fd_sc_hd__buf_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15262_ _08688_/X _15262_/D VGND VGND VPWR VPWR _15262_/Q sky130_fd_sc_hd__dfxtp_1
X_12474_ _12509_/A VGND VGND VPWR VPWR _12480_/B sky130_fd_sc_hd__clkbuf_4
X_14213_ _14666_/Q _15242_/Q _14730_/Q _14698_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14213_/X sky130_fd_sc_hd__mux4_2
X_11425_ _11436_/A VGND VGND VPWR VPWR _11425_/X sky130_fd_sc_hd__clkbuf_1
X_15193_ _08962_/X _15193_/D VGND VGND VPWR VPWR _15193_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_7 data_address[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14144_ _15185_/Q _15153_/Q _14769_/Q _14801_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14144_/X sky130_fd_sc_hd__mux4_1
X_11356_ _14585_/Q _11354_/X _11108_/X _11355_/X VGND VGND VPWR VPWR _14585_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10307_ _10319_/A VGND VGND VPWR VPWR _10307_/X sky130_fd_sc_hd__clkbuf_1
X_14075_ _15128_/Q _15352_/Q _15320_/Q _15288_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14075_/X sky130_fd_sc_hd__mux4_1
X_11287_ _14605_/Q _11284_/X _11161_/X _11286_/X VGND VGND VPWR VPWR _14605_/D sky130_fd_sc_hd__a22o_1
XFILLER_140_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13026_ _15669_/Q _07642_/A _12556_/A _07909_/C _07184_/X VGND VGND VPWR VPWR _15669_/D
+ sky130_fd_sc_hd__o221a_1
X_10238_ _10248_/A VGND VGND VPWR VPWR _10238_/X sky130_fd_sc_hd__buf_1
XFILLER_67_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10169_ _10171_/A VGND VGND VPWR VPWR _10169_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14977_ _09818_/X _14977_/D VGND VGND VPWR VPWR _14977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13928_ _14503_/Q _14471_/Q _14439_/Q _14407_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13928_/X sky130_fd_sc_hd__mux4_2
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13859_ _14830_/Q _14862_/Q _14894_/Q _14926_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13859_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07380_ _07510_/B _07322_/X _12569_/A _07373_/X VGND VGND VPWR VPWR _07380_/X sky130_fd_sc_hd__o22a_1
X_15529_ _15579_/CLK _15529_/D VGND VGND VPWR VPWR _15529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09050_ _15168_/Q _09041_/X _08793_/X _09044_/X VGND VGND VPWR VPWR _15168_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08001_ _08049_/A VGND VGND VPWR VPWR _08032_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09952_ _09952_/A VGND VGND VPWR VPWR _09961_/A sky130_fd_sc_hd__buf_1
XFILLER_104_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08903_ _08908_/A VGND VGND VPWR VPWR _08903_/X sky130_fd_sc_hd__clkbuf_1
X_09883_ _09885_/A VGND VGND VPWR VPWR _09883_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08834_ _09206_/A VGND VGND VPWR VPWR _08834_/X sky130_fd_sc_hd__buf_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08765_ _08765_/A VGND VGND VPWR VPWR _08770_/A sky130_fd_sc_hd__buf_1
X_07716_ _07715_/X _13140_/X _07715_/X _13140_/X VGND VGND VPWR VPWR _07871_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_26_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08696_ _08705_/A VGND VGND VPWR VPWR _08701_/A sky130_fd_sc_hd__buf_1
X_07647_ _07647_/A VGND VGND VPWR VPWR _07687_/A sky130_fd_sc_hd__buf_1
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07578_ _07582_/A VGND VGND VPWR VPWR _07581_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09317_ _15102_/Q _09311_/X _09176_/X _09314_/X VGND VGND VPWR VPWR _15102_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09248_ _09248_/A VGND VGND VPWR VPWR _09274_/A sky130_fd_sc_hd__buf_1
XFILLER_107_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09179_ _09187_/A VGND VGND VPWR VPWR _09179_/X sky130_fd_sc_hd__buf_1
XFILLER_135_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11210_ _11210_/A VGND VGND VPWR VPWR _11210_/X sky130_fd_sc_hd__buf_1
X_12190_ _12190_/A _12190_/B VGND VGND VPWR VPWR _12750_/A sky130_fd_sc_hd__or2_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11141_ _11216_/A VGND VGND VPWR VPWR _11168_/A sky130_fd_sc_hd__buf_2
XFILLER_1_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11072_ _14657_/Q _11064_/X _11071_/X _11068_/X VGND VGND VPWR VPWR _14657_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14900_ _10123_/X _14900_/D VGND VGND VPWR VPWR _14900_/Q sky130_fd_sc_hd__dfxtp_1
X_10023_ _10023_/A VGND VGND VPWR VPWR _10050_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14831_ _10382_/X _14831_/D VGND VGND VPWR VPWR _14831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14762_ _10636_/X _14762_/D VGND VGND VPWR VPWR _14762_/Q sky130_fd_sc_hd__dfxtp_1
X_11974_ _11994_/A VGND VGND VPWR VPWR _11981_/A sky130_fd_sc_hd__buf_1
XFILLER_17_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13713_ _14684_/Q _15260_/Q _14748_/Q _14716_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13713_/X sky130_fd_sc_hd__mux4_1
X_10925_ _10937_/A VGND VGND VPWR VPWR _10925_/X sky130_fd_sc_hd__buf_1
X_14693_ _10941_/X _14693_/D VGND VGND VPWR VPWR _14693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13644_ _14276_/X _14281_/X _13648_/S VGND VGND VPWR VPWR _13644_/X sky130_fd_sc_hd__mux2_1
X_10856_ _10875_/A VGND VGND VPWR VPWR _10856_/X sky130_fd_sc_hd__buf_1
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _13574_/X _13078_/X _14337_/Q VGND VGND VPWR VPWR _13575_/X sky130_fd_sc_hd__mux2_1
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10787_ _10787_/A VGND VGND VPWR VPWR _11533_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15314_ _08451_/X _15314_/D VGND VGND VPWR VPWR _15314_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12526_ _15560_/Q VGND VGND VPWR VPWR _12962_/B sky130_fd_sc_hd__clkbuf_2
X_15245_ _08740_/X _15245_/D VGND VGND VPWR VPWR _15245_/Q sky130_fd_sc_hd__dfxtp_1
X_12457_ _12874_/A VGND VGND VPWR VPWR _12819_/A sky130_fd_sc_hd__buf_1
XFILLER_8_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11408_ _11424_/A VGND VGND VPWR VPWR _11413_/A sky130_fd_sc_hd__buf_1
XFILLER_126_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15176_ _09021_/X _15176_/D VGND VGND VPWR VPWR _15176_/Q sky130_fd_sc_hd__dfxtp_1
X_12388_ _12392_/A VGND VGND VPWR VPWR _12388_/X sky130_fd_sc_hd__buf_4
X_14127_ _14643_/Q _14611_/Q _14579_/Q _15379_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14127_/X sky130_fd_sc_hd__mux4_2
XFILLER_125_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11339_ _14590_/Q _11332_/X _11087_/X _11335_/X VGND VGND VPWR VPWR _14590_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14058_ _14522_/Q _14490_/Q _14458_/Q _14426_/Q _14395_/Q _14060_/S1 VGND VGND VPWR
+ VPWR _14058_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13009_ _14353_/Q VGND VGND VPWR VPWR _13009_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_opt_4_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR clkbuf_opt_4_clk/X sky130_fd_sc_hd__clkbuf_16
X_08550_ _09296_/A _08550_/B VGND VGND VPWR VPWR _08563_/A sky130_fd_sc_hd__or2_2
X_07501_ _07613_/A VGND VGND VPWR VPWR _07511_/A sky130_fd_sc_hd__buf_1
XFILLER_51_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08481_ _08481_/A VGND VGND VPWR VPWR _08520_/A sky130_fd_sc_hd__buf_1
XFILLER_90_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07432_ _07432_/A _13627_/X VGND VGND VPWR VPWR _15567_/D sky130_fd_sc_hd__and2_1
XFILLER_90_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07363_ _07363_/A VGND VGND VPWR VPWR _07363_/X sky130_fd_sc_hd__buf_1
X_09102_ _15154_/Q _09095_/X _08856_/X _09096_/X VGND VGND VPWR VPWR _15154_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07294_ _14375_/Q VGND VGND VPWR VPWR _07559_/A sky130_fd_sc_hd__inv_2
XFILLER_136_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09033_ _09059_/A VGND VGND VPWR VPWR _09038_/A sky130_fd_sc_hd__buf_1
XFILLER_117_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09935_ _14945_/Q _09927_/X _09934_/X _09931_/X VGND VGND VPWR VPWR _14945_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09866_ _14964_/Q _09856_/X _09607_/X _09858_/X VGND VGND VPWR VPWR _14964_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08817_ _09188_/A VGND VGND VPWR VPWR _08817_/X sky130_fd_sc_hd__buf_1
XFILLER_100_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09797_ _09797_/A VGND VGND VPWR VPWR _09797_/X sky130_fd_sc_hd__buf_1
XFILLER_27_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08748_ _08752_/A VGND VGND VPWR VPWR _08748_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_205 _13516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_216 _13019_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_227 _08741_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_238 _11239_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08679_ _08702_/A VGND VGND VPWR VPWR _08679_/X sky130_fd_sc_hd__buf_1
XANTENNA_249 _11951_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10710_ _10725_/A VGND VGND VPWR VPWR _10721_/A sky130_fd_sc_hd__buf_1
XFILLER_41_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11690_ _11703_/A VGND VGND VPWR VPWR _11691_/A sky130_fd_sc_hd__buf_1
X_10641_ _10645_/A VGND VGND VPWR VPWR _10641_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13360_ _13359_/X _13361_/X _15565_/Q VGND VGND VPWR VPWR _13360_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10572_ _10574_/A VGND VGND VPWR VPWR _10572_/X sky130_fd_sc_hd__clkbuf_1
X_12311_ _12681_/A VGND VGND VPWR VPWR _12663_/A sky130_fd_sc_hd__buf_1
XFILLER_6_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13291_ _13290_/X _13292_/X _15565_/Q VGND VGND VPWR VPWR _13291_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15030_ _09591_/X _15030_/D VGND VGND VPWR VPWR _15030_/Q sky130_fd_sc_hd__dfxtp_1
X_12242_ _12246_/A VGND VGND VPWR VPWR _12820_/A sky130_fd_sc_hd__buf_1
XFILLER_5_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12173_ _15574_/Q VGND VGND VPWR VPWR _12726_/A sky130_fd_sc_hd__inv_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11124_ _14646_/Q _11120_/X _11121_/X _11123_/X VGND VGND VPWR VPWR _14646_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11055_ _14660_/Q _10951_/A _10828_/X _10954_/A VGND VGND VPWR VPWR _14660_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10006_ _10032_/A VGND VGND VPWR VPWR _10015_/A sky130_fd_sc_hd__buf_1
XFILLER_92_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14814_ _10458_/X _14814_/D VGND VGND VPWR VPWR _14814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14745_ _10715_/X _14745_/D VGND VGND VPWR VPWR _14745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11957_ _11987_/A VGND VGND VPWR VPWR _11977_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10908_ _14703_/Q _10904_/X _10771_/X _10905_/X VGND VGND VPWR VPWR _14703_/D sky130_fd_sc_hd__a22o_1
X_14676_ _11003_/X _14676_/D VGND VGND VPWR VPWR _14676_/Q sky130_fd_sc_hd__dfxtp_1
X_11888_ _14442_/Q _11886_/X _08064_/A _11887_/X VGND VGND VPWR VPWR _14442_/D sky130_fd_sc_hd__a22o_1
X_13627_ _13626_/X _13065_/X _14337_/Q VGND VGND VPWR VPWR _13627_/X sky130_fd_sc_hd__mux2_1
Xrepeater30 _13945_/S0 VGND VGND VPWR VPWR _13919_/S0 sky130_fd_sc_hd__clkbuf_16
XFILLER_20_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater41 _14210_/S1 VGND VGND VPWR VPWR _14238_/S1 sky130_fd_sc_hd__clkbuf_16
X_10839_ _10851_/A VGND VGND VPWR VPWR _10840_/A sky130_fd_sc_hd__buf_1
Xrepeater52 _14395_/Q VGND VGND VPWR VPWR _14055_/S0 sky130_fd_sc_hd__buf_12
X_13558_ _13557_/X _14327_/D _15506_/Q VGND VGND VPWR VPWR _13558_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12509_ _12509_/A _12509_/B VGND VGND VPWR VPWR _12509_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13489_ _13488_/X rdata[11] _13516_/S VGND VGND VPWR VPWR _13489_/X sky130_fd_sc_hd__mux2_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15228_ _08811_/X _15228_/D VGND VGND VPWR VPWR _15228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15159_ _09081_/X _15159_/D VGND VGND VPWR VPWR _15159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07981_ _07981_/A VGND VGND VPWR VPWR _07981_/X sky130_fd_sc_hd__buf_1
XFILLER_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09720_ _09722_/A VGND VGND VPWR VPWR _09720_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09651_ _09964_/A VGND VGND VPWR VPWR _09860_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_68_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08602_ _15285_/Q _08597_/X _08434_/X _08599_/X VGND VGND VPWR VPWR _15285_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09582_ _09582_/A VGND VGND VPWR VPWR _09582_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08533_ _14306_/Q VGND VGND VPWR VPWR _10823_/A sky130_fd_sc_hd__buf_1
XFILLER_70_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ _14317_/Q VGND VGND VPWR VPWR _10765_/A sky130_fd_sc_hd__buf_1
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07415_ _07415_/A _13579_/X VGND VGND VPWR VPWR _15579_/D sky130_fd_sc_hd__and2_1
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ _10707_/A VGND VGND VPWR VPWR _09188_/A sky130_fd_sc_hd__buf_1
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07346_ _14389_/Q VGND VGND VPWR VPWR _07497_/B sky130_fd_sc_hd__inv_2
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07277_ _07278_/A _07277_/B VGND VGND VPWR VPWR _15617_/D sky130_fd_sc_hd__nor2_1
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09016_ _09025_/A VGND VGND VPWR VPWR _09016_/X sky130_fd_sc_hd__buf_1
XFILLER_152_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09918_ _09952_/A VGND VGND VPWR VPWR _09933_/A sky130_fd_sc_hd__buf_1
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09849_ _09849_/A VGND VGND VPWR VPWR _09854_/A sky130_fd_sc_hd__buf_1
XFILLER_58_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12860_ _12860_/A _12860_/B VGND VGND VPWR VPWR _12861_/A sky130_fd_sc_hd__or2_1
X_11811_ _11811_/A VGND VGND VPWR VPWR _11874_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12791_ _12791_/A VGND VGND VPWR VPWR _12791_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14530_ _11573_/X _14530_/D VGND VGND VPWR VPWR _14530_/Q sky130_fd_sc_hd__dfxtp_1
X_11742_ _11742_/A VGND VGND VPWR VPWR _11742_/X sky130_fd_sc_hd__clkbuf_1
X_14461_ _11822_/X _14461_/D VGND VGND VPWR VPWR _14461_/Q sky130_fd_sc_hd__dfxtp_1
X_11673_ _11673_/A VGND VGND VPWR VPWR _11673_/X sky130_fd_sc_hd__buf_1
X_13412_ _13414_/X _13413_/X _13415_/S VGND VGND VPWR VPWR _13412_/X sky130_fd_sc_hd__mux2_1
X_10624_ _14766_/Q _10616_/X _10389_/X _10617_/X VGND VGND VPWR VPWR _14766_/D sky130_fd_sc_hd__a22o_1
X_14392_ _14392_/CLK instruction[29] VGND VGND VPWR VPWR _14392_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13343_ _13342_/X _13344_/X _15565_/Q VGND VGND VPWR VPWR _13343_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10555_ _10555_/A VGND VGND VPWR VPWR _10578_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13274_ _13275_/X _12883_/B _15564_/Q VGND VGND VPWR VPWR _13274_/X sky130_fd_sc_hd__mux2_2
X_10486_ _10506_/A VGND VGND VPWR VPWR _10486_/X sky130_fd_sc_hd__buf_1
XFILLER_142_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15013_ _09685_/X _15013_/D VGND VGND VPWR VPWR _15013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12225_ _15562_/Q _12157_/X _12815_/A _12106_/A VGND VGND VPWR VPWR _12225_/X sky130_fd_sc_hd__o22a_1
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12156_ _12156_/A VGND VGND VPWR VPWR _12157_/A sky130_fd_sc_hd__buf_1
XFILLER_111_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11107_ _11107_/A VGND VGND VPWR VPWR _11107_/X sky130_fd_sc_hd__buf_1
XFILLER_96_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12087_ _15552_/Q _12087_/B VGND VGND VPWR VPWR _12087_/Y sky130_fd_sc_hd__nor2_2
XFILLER_96_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11038_ _11047_/A VGND VGND VPWR VPWR _11038_/X sky130_fd_sc_hd__buf_1
XFILLER_65_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12989_ _15514_/Q _12568_/A _15517_/Q _07366_/A VGND VGND VPWR VPWR _12989_/X sky130_fd_sc_hd__o22a_1
XFILLER_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14728_ _10807_/X _14728_/D VGND VGND VPWR VPWR _14728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14659_ _11058_/X _14659_/D VGND VGND VPWR VPWR _14659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07200_ _07235_/A VGND VGND VPWR VPWR _07200_/X sky130_fd_sc_hd__buf_2
X_08180_ _08180_/A VGND VGND VPWR VPWR _08189_/A sky130_fd_sc_hd__buf_1
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07131_ _13113_/X VGND VGND VPWR VPWR _07259_/B sky130_fd_sc_hd__inv_2
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07964_ _15421_/Q _07949_/X _07963_/X _07954_/X VGND VGND VPWR VPWR _15421_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09703_ _09713_/A VGND VGND VPWR VPWR _09716_/A sky130_fd_sc_hd__inv_2
XFILLER_28_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07895_ _07895_/A _07895_/B VGND VGND VPWR VPWR _07895_/X sky130_fd_sc_hd__or2_1
XFILLER_55_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09634_ _09634_/A VGND VGND VPWR VPWR _09647_/A sky130_fd_sc_hd__buf_1
XFILLER_83_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09565_ _09580_/A VGND VGND VPWR VPWR _09565_/X sky130_fd_sc_hd__buf_1
XFILLER_24_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08516_ _10808_/A VGND VGND VPWR VPWR _09271_/A sky130_fd_sc_hd__buf_1
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09496_ _09505_/A VGND VGND VPWR VPWR _09496_/X sky130_fd_sc_hd__buf_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08447_ _10750_/A VGND VGND VPWR VPWR _09224_/A sky130_fd_sc_hd__buf_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08378_ _15326_/Q _08366_/X _08377_/X _08372_/X VGND VGND VPWR VPWR _15326_/D sky130_fd_sc_hd__a22o_1
X_07329_ _07337_/A _07329_/B VGND VGND VPWR VPWR _15603_/D sky130_fd_sc_hd__nor2_1
XFILLER_136_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10340_ _10340_/A VGND VGND VPWR VPWR _10340_/X sky130_fd_sc_hd__buf_1
XFILLER_125_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10271_ _10931_/A VGND VGND VPWR VPWR _10492_/A sky130_fd_sc_hd__buf_1
XFILLER_151_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12010_ _12010_/A VGND VGND VPWR VPWR _12010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13961_ _13957_/X _13958_/X _13959_/X _13960_/X _07533_/A _14402_/Q VGND VGND VPWR
+ VPWR _13961_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12912_ _12724_/X _12172_/X _12725_/A _12726_/A VGND VGND VPWR VPWR _12914_/C sky130_fd_sc_hd__o22a_1
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13892_ _15210_/Q _14538_/Q _14986_/Q _15402_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13892_/X sky130_fd_sc_hd__mux4_2
XFILLER_47_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15631_ _15663_/CLK _15631_/D VGND VGND VPWR VPWR pc[26] sky130_fd_sc_hd__dfxtp_4
X_12843_ _12843_/A VGND VGND VPWR VPWR _12847_/B sky130_fd_sc_hd__buf_1
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15562_ _15578_/CLK _15562_/D VGND VGND VPWR VPWR _15562_/Q sky130_fd_sc_hd__dfxtp_4
X_12774_ _12774_/A VGND VGND VPWR VPWR _12775_/A sky130_fd_sc_hd__buf_1
XFILLER_61_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14513_ _11638_/X _14513_/D VGND VGND VPWR VPWR _14513_/Q sky130_fd_sc_hd__dfxtp_1
X_11725_ _11725_/A VGND VGND VPWR VPWR _11746_/A sky130_fd_sc_hd__clkbuf_2
X_15493_ _15579_/CLK _15493_/D VGND VGND VPWR VPWR wdata[19] sky130_fd_sc_hd__dfxtp_4
XFILLER_70_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14444_ _11879_/X _14444_/D VGND VGND VPWR VPWR _14444_/Q sky130_fd_sc_hd__dfxtp_1
X_11656_ _11658_/A VGND VGND VPWR VPWR _11656_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10607_ _10616_/A VGND VGND VPWR VPWR _10607_/X sky130_fd_sc_hd__buf_1
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14375_ _14375_/CLK instruction[4] VGND VGND VPWR VPWR _14375_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ _11587_/A VGND VGND VPWR VPWR _11598_/A sky130_fd_sc_hd__buf_1
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13326_ _13325_/X _13334_/X _13393_/S VGND VGND VPWR VPWR _13326_/X sky130_fd_sc_hd__mux2_1
X_10538_ _10540_/A VGND VGND VPWR VPWR _10538_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13257_ _13258_/X _13282_/X _13408_/S VGND VGND VPWR VPWR _13257_/X sky130_fd_sc_hd__mux2_1
X_10469_ _14811_/Q _10465_/X _10332_/X _10466_/X VGND VGND VPWR VPWR _14811_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12208_ _12773_/A _12275_/B _12207_/Y VGND VGND VPWR VPWR _12746_/A sky130_fd_sc_hd__a21oi_1
X_13188_ _13191_/X _13211_/X _15563_/Q VGND VGND VPWR VPWR _13188_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12139_ _15578_/Q VGND VGND VPWR VPWR _12139_/X sky130_fd_sc_hd__buf_1
XFILLER_69_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07680_ _07680_/A VGND VGND VPWR VPWR _07706_/A sky130_fd_sc_hd__buf_1
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09350_ _15093_/Q _09345_/X _09216_/X _09347_/X VGND VGND VPWR VPWR _15093_/D sky130_fd_sc_hd__a22o_1
X_08301_ _15343_/Q _08291_/X _08036_/X _08292_/X VGND VGND VPWR VPWR _15343_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09281_ _09281_/A VGND VGND VPWR VPWR _09307_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08232_ _08264_/A VGND VGND VPWR VPWR _08255_/A sky130_fd_sc_hd__clkbuf_4
X_08163_ _08169_/A VGND VGND VPWR VPWR _08163_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07114_ _07642_/A _15668_/Q _07909_/C data_address[0] _07291_/A VGND VGND VPWR VPWR
+ _15668_/D sky130_fd_sc_hd__o221a_1
X_08094_ _14305_/Q VGND VGND VPWR VPWR _08095_/A sky130_fd_sc_hd__buf_1
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08996_ _08998_/A VGND VGND VPWR VPWR _08996_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07947_ _07947_/A VGND VGND VPWR VPWR _08045_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07878_ _07878_/A _07878_/B VGND VGND VPWR VPWR _07878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09617_ _10371_/A VGND VGND VPWR VPWR _09617_/X sky130_fd_sc_hd__buf_1
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09548_ _09644_/A VGND VGND VPWR VPWR _09580_/A sky130_fd_sc_hd__buf_2
XFILLER_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ _09499_/A VGND VGND VPWR VPWR _09484_/A sky130_fd_sc_hd__buf_2
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11510_ _11510_/A VGND VGND VPWR VPWR _11510_/X sky130_fd_sc_hd__buf_1
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12490_ _15559_/Q VGND VGND VPWR VPWR _12491_/A sky130_fd_sc_hd__inv_2
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ _11469_/A VGND VGND VPWR VPWR _11454_/A sky130_fd_sc_hd__buf_1
XFILLER_149_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14160_ _14960_/Q _15056_/Q _15024_/Q _15088_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14160_/X sky130_fd_sc_hd__mux4_2
XFILLER_109_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11372_ _14580_/Q _11364_/X _11130_/X _11366_/X VGND VGND VPWR VPWR _14580_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13111_ _15657_/Q data_address[22] _15667_/Q VGND VGND VPWR VPWR _13111_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10323_ _10331_/A VGND VGND VPWR VPWR _10323_/X sky130_fd_sc_hd__clkbuf_1
X_14091_ _14087_/X _14088_/X _14089_/X _14090_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14091_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13042_ wdata[15] rdata[15] ren VGND VGND VPWR VPWR _14319_/D sky130_fd_sc_hd__mux2_1
X_10254_ _14862_/Q _10247_/X _10020_/X _10248_/X VGND VGND VPWR VPWR _14862_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10185_ _10197_/A VGND VGND VPWR VPWR _10186_/A sky130_fd_sc_hd__buf_1
XFILLER_78_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14993_ _09761_/X _14993_/D VGND VGND VPWR VPWR _14993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13944_ _15173_/Q _15141_/Q _14757_/Q _14789_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13944_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13875_ _15116_/Q _15340_/Q _15308_/Q _15276_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13875_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12826_ _12826_/A VGND VGND VPWR VPWR _12826_/X sky130_fd_sc_hd__buf_1
X_15614_ _15646_/CLK _15614_/D VGND VGND VPWR VPWR pc[9] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12757_ _12752_/X _12179_/X _12753_/X _12756_/X VGND VGND VPWR VPWR _12757_/Y sky130_fd_sc_hd__o22ai_1
X_15545_ _15578_/CLK _15545_/D VGND VGND VPWR VPWR _15545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11708_ _11712_/A VGND VGND VPWR VPWR _11708_/X sky130_fd_sc_hd__clkbuf_1
X_15476_ _15521_/CLK _15476_/D VGND VGND VPWR VPWR wdata[2] sky130_fd_sc_hd__dfxtp_2
X_12688_ _12684_/X _12735_/A _12735_/B _12273_/A VGND VGND VPWR VPWR _12689_/B sky130_fd_sc_hd__a31o_1
XFILLER_129_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14427_ _11939_/X _14427_/D VGND VGND VPWR VPWR _14427_/Q sky130_fd_sc_hd__dfxtp_1
X_11639_ _14513_/Q _11633_/X _11510_/X _11634_/X VGND VGND VPWR VPWR _14513_/D sky130_fd_sc_hd__a22o_1
XFILLER_128_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358_ _15654_/CLK pc[19] VGND VGND VPWR VPWR _14358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13309_ _13308_/X _13310_/X _15565_/Q VGND VGND VPWR VPWR _13309_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14289_ _14819_/Q _14851_/Q _14883_/Q _14915_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14289_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08850_ _08855_/A VGND VGND VPWR VPWR _08850_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07801_ _07668_/A _07800_/Y _07668_/Y _07800_/A _07640_/A VGND VGND VPWR VPWR _15456_/D
+ sky130_fd_sc_hd__o221a_1
X_08781_ _08796_/A VGND VGND VPWR VPWR _08782_/A sky130_fd_sc_hd__buf_1
XFILLER_111_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07732_ _13143_/X _07728_/B _07728_/Y _07731_/X VGND VGND VPWR VPWR _07733_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07663_ _07663_/A VGND VGND VPWR VPWR _07663_/X sky130_fd_sc_hd__clkbuf_1
X_09402_ _09402_/A VGND VGND VPWR VPWR _09407_/A sky130_fd_sc_hd__buf_1
X_07594_ _07595_/A _13072_/X VGND VGND VPWR VPWR _15487_/D sky130_fd_sc_hd__and2_1
XFILLER_34_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09333_ _09342_/A VGND VGND VPWR VPWR _09340_/A sky130_fd_sc_hd__buf_1
XFILLER_34_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09264_ _09276_/A VGND VGND VPWR VPWR _09264_/X sky130_fd_sc_hd__buf_1
X_08215_ _15363_/Q _08109_/A _08099_/X _08112_/A VGND VGND VPWR VPWR _15363_/D sky130_fd_sc_hd__a22o_1
X_09195_ _09195_/A VGND VGND VPWR VPWR _09195_/X sky130_fd_sc_hd__buf_1
XFILLER_147_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08146_ _08148_/A VGND VGND VPWR VPWR _08146_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08077_ _08077_/A VGND VGND VPWR VPWR _08077_/X sky130_fd_sc_hd__buf_1
XFILLER_105_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08979_ _15189_/Q _08974_/X _08844_/X _08976_/X VGND VGND VPWR VPWR _15189_/D sky130_fd_sc_hd__a22o_1
XFILLER_76_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11990_ _11992_/A VGND VGND VPWR VPWR _11990_/X sky130_fd_sc_hd__clkbuf_1
X_10941_ _10941_/A VGND VGND VPWR VPWR _10941_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13660_ _14978_/Q _15074_/Q _15042_/Q _15106_/Q _13740_/S0 _07541_/A VGND VGND VPWR
+ VPWR _13660_/X sky130_fd_sc_hd__mux4_2
X_10872_ _10892_/A VGND VGND VPWR VPWR _10879_/A sky130_fd_sc_hd__buf_1
XFILLER_25_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12611_ _12611_/A VGND VGND VPWR VPWR _12611_/X sky130_fd_sc_hd__clkbuf_4
X_13591_ _13590_/X _13074_/X _14337_/Q VGND VGND VPWR VPWR _13591_/X sky130_fd_sc_hd__mux2_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15330_ _08339_/X _15330_/D VGND VGND VPWR VPWR _15330_/Q sky130_fd_sc_hd__dfxtp_1
X_12542_ _15471_/Q VGND VGND VPWR VPWR _12545_/A sky130_fd_sc_hd__inv_2
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15261_ _08690_/X _15261_/D VGND VGND VPWR VPWR _15261_/Q sky130_fd_sc_hd__dfxtp_1
X_12473_ _12473_/A VGND VGND VPWR VPWR _12480_/A sky130_fd_sc_hd__buf_1
XFILLER_8_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14212_ _15210_/Q _14538_/Q _14986_/Q _15402_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14212_/X sky130_fd_sc_hd__mux4_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11424_ _11424_/A VGND VGND VPWR VPWR _11436_/A sky130_fd_sc_hd__clkbuf_2
X_15192_ _08966_/X _15192_/D VGND VGND VPWR VPWR _15192_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_8 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14143_ _14673_/Q _15249_/Q _14737_/Q _14705_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14143_/X sky130_fd_sc_hd__mux4_2
X_11355_ _11355_/A VGND VGND VPWR VPWR _11355_/X sky130_fd_sc_hd__buf_1
XFILLER_153_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10306_ _10334_/A VGND VGND VPWR VPWR _10319_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14074_ _15192_/Q _15160_/Q _14776_/Q _14808_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14074_/X sky130_fd_sc_hd__mux4_2
X_11286_ _11304_/A VGND VGND VPWR VPWR _11286_/X sky130_fd_sc_hd__buf_1
XFILLER_140_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13025_ _14369_/Q VGND VGND VPWR VPWR _13025_/Y sky130_fd_sc_hd__inv_2
X_10237_ _10247_/A VGND VGND VPWR VPWR _10237_/X sky130_fd_sc_hd__buf_1
XFILLER_140_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10168_ _14887_/Q _10166_/X _10051_/X _10167_/X VGND VGND VPWR VPWR _14887_/D sky130_fd_sc_hd__a22o_1
XFILLER_120_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14976_ _09820_/X _14976_/D VGND VGND VPWR VPWR _14976_/Q sky130_fd_sc_hd__dfxtp_1
X_10099_ _14908_/Q _10097_/X _09958_/X _10098_/X VGND VGND VPWR VPWR _14908_/D sky130_fd_sc_hd__a22o_1
XFILLER_47_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13927_ _14631_/Q _14599_/Q _14567_/Q _15367_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13927_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13858_ _14510_/Q _14478_/Q _14446_/Q _14414_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13858_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12809_ _12805_/X _12235_/X _12753_/X _12808_/X VGND VGND VPWR VPWR _12809_/Y sky130_fd_sc_hd__o22ai_1
X_13789_ _14837_/Q _14869_/Q _14901_/Q _14933_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13789_/X sky130_fd_sc_hd__mux4_2
XFILLER_50_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15528_ _15599_/CLK _15528_/D VGND VGND VPWR VPWR _15528_/Q sky130_fd_sc_hd__dfxtp_1
X_15459_ _15604_/CLK _15459_/D VGND VGND VPWR VPWR _15459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08000_ _08000_/A VGND VGND VPWR VPWR _08000_/X sky130_fd_sc_hd__buf_1
XFILLER_128_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09951_ _14942_/Q _09943_/X _09950_/X _09947_/X VGND VGND VPWR VPWR _14942_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08902_ _15208_/Q _08890_/X _08901_/X _08892_/X VGND VGND VPWR VPWR _15208_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09882_ _14959_/Q _09877_/X _09632_/X _09878_/X VGND VGND VPWR VPWR _14959_/D sky130_fd_sc_hd__a22o_1
X_08833_ _08843_/A VGND VGND VPWR VPWR _08833_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08764_ _15239_/Q _08762_/X _08523_/X _08763_/X VGND VGND VPWR VPWR _15239_/D sky130_fd_sc_hd__a22o_1
X_07715_ _07715_/A VGND VGND VPWR VPWR _07715_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08695_ _15260_/Q _08693_/X _08390_/X _08694_/X VGND VGND VPWR VPWR _15260_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07646_ _07679_/A VGND VGND VPWR VPWR _07647_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_80_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07577_ _07577_/A _13083_/X VGND VGND VPWR VPWR _15498_/D sky130_fd_sc_hd__and2_1
XFILLER_80_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09316_ _09318_/A VGND VGND VPWR VPWR _09316_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09247_ _09254_/A VGND VGND VPWR VPWR _09247_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09178_ _09190_/A VGND VGND VPWR VPWR _09187_/A sky130_fd_sc_hd__buf_1
XFILLER_147_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08129_ _08129_/A VGND VGND VPWR VPWR _08129_/X sky130_fd_sc_hd__clkbuf_1
X_11140_ _11140_/A VGND VGND VPWR VPWR _11216_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11071_ _11437_/A VGND VGND VPWR VPWR _11071_/X sky130_fd_sc_hd__buf_1
XFILLER_89_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10022_ _10029_/A VGND VGND VPWR VPWR _10022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14830_ _10388_/X _14830_/D VGND VGND VPWR VPWR _14830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11973_ _11973_/A VGND VGND VPWR VPWR _11994_/A sky130_fd_sc_hd__clkbuf_4
X_14761_ _10641_/X _14761_/D VGND VGND VPWR VPWR _14761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10924_ _10936_/A VGND VGND VPWR VPWR _10924_/X sky130_fd_sc_hd__buf_1
X_13712_ _15228_/Q _14556_/Q _15004_/Q _15420_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13712_/X sky130_fd_sc_hd__mux4_1
X_14692_ _10944_/X _14692_/D VGND VGND VPWR VPWR _14692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10855_ _10915_/A VGND VGND VPWR VPWR _10875_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13643_ _13642_/X _13061_/X _14337_/Q VGND VGND VPWR VPWR _13643_/X sky130_fd_sc_hd__mux2_1
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13574_ _13573_/X _14323_/D _15506_/Q VGND VGND VPWR VPWR _13574_/X sky130_fd_sc_hd__mux2_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10786_ _10786_/A VGND VGND VPWR VPWR _10786_/X sky130_fd_sc_hd__clkbuf_1
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12525_ _12962_/A _12522_/X _12336_/X _12496_/X _12521_/X VGND VGND VPWR VPWR _12525_/X
+ sky130_fd_sc_hd__o32a_1
X_15313_ _08457_/X _15313_/D VGND VGND VPWR VPWR _15313_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12456_ _12456_/A VGND VGND VPWR VPWR _12846_/B sky130_fd_sc_hd__buf_1
X_15244_ _08748_/X _15244_/D VGND VGND VPWR VPWR _15244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11407_ _11407_/A VGND VGND VPWR VPWR _11424_/A sky130_fd_sc_hd__buf_1
X_15175_ _09024_/X _15175_/D VGND VGND VPWR VPWR _15175_/Q sky130_fd_sc_hd__dfxtp_1
X_12387_ _15555_/Q VGND VGND VPWR VPWR _12392_/A sky130_fd_sc_hd__inv_2
X_14126_ _14122_/X _14123_/X _14124_/X _14125_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14126_/X sky130_fd_sc_hd__mux4_2
X_11338_ _11342_/A VGND VGND VPWR VPWR _11338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14057_ _14650_/Q _14618_/Q _14586_/Q _15386_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14057_/X sky130_fd_sc_hd__mux4_2
X_11269_ _11269_/A VGND VGND VPWR VPWR _11269_/X sky130_fd_sc_hd__clkbuf_1
X_13008_ _14352_/Q VGND VGND VPWR VPWR _13008_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14959_ _09881_/X _14959_/D VGND VGND VPWR VPWR _14959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07500_ _07500_/A _12563_/C VGND VGND VPWR VPWR _15521_/D sky130_fd_sc_hd__nor2_1
X_08480_ _08489_/A VGND VGND VPWR VPWR _08480_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07431_ _07432_/A _13623_/X VGND VGND VPWR VPWR _15568_/D sky130_fd_sc_hd__and2_1
X_07362_ _07377_/A _07362_/B VGND VGND VPWR VPWR _15597_/D sky130_fd_sc_hd__nor2_1
X_09101_ _09105_/A VGND VGND VPWR VPWR _09101_/X sky130_fd_sc_hd__clkbuf_1
X_07293_ _14377_/Q VGND VGND VPWR VPWR _07559_/C sky130_fd_sc_hd__buf_1
XFILLER_149_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09032_ _09068_/A VGND VGND VPWR VPWR _09059_/A sky130_fd_sc_hd__buf_2
XFILLER_117_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09934_ _10303_/A VGND VGND VPWR VPWR _09934_/X sky130_fd_sc_hd__buf_1
XFILLER_104_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09865_ _09867_/A VGND VGND VPWR VPWR _09865_/X sky130_fd_sc_hd__clkbuf_1
X_08816_ _08816_/A VGND VGND VPWR VPWR _08816_/X sky130_fd_sc_hd__clkbuf_1
X_09796_ _09802_/A VGND VGND VPWR VPWR _09796_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08747_ _08765_/A VGND VGND VPWR VPWR _08752_/A sky130_fd_sc_hd__buf_1
XANTENNA_206 _13512_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_217 _13021_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_228 _08743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08678_ _08741_/A VGND VGND VPWR VPWR _08702_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_239 _11337_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07629_ _07630_/A _07629_/B VGND VGND VPWR VPWR _15469_/D sky130_fd_sc_hd__nor2_1
XFILLER_81_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10640_ _10640_/A VGND VGND VPWR VPWR _10645_/A sky130_fd_sc_hd__buf_1
XFILLER_139_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10571_ _14782_/Q _10564_/X _10320_/X _10567_/X VGND VGND VPWR VPWR _14782_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12310_ _12426_/A VGND VGND VPWR VPWR _12681_/A sky130_fd_sc_hd__buf_1
X_13290_ _13289_/X _13294_/X _13393_/S VGND VGND VPWR VPWR _13290_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12241_ _15535_/Q VGND VGND VPWR VPWR _12246_/A sky130_fd_sc_hd__inv_2
XFILLER_5_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12172_ _15574_/Q VGND VGND VPWR VPWR _12172_/X sky130_fd_sc_hd__buf_1
X_11123_ _11149_/A VGND VGND VPWR VPWR _11123_/X sky130_fd_sc_hd__buf_1
XFILLER_1_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11054_ _11054_/A VGND VGND VPWR VPWR _11054_/X sky130_fd_sc_hd__buf_1
XFILLER_77_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10005_ _10044_/A VGND VGND VPWR VPWR _10032_/A sky130_fd_sc_hd__buf_2
XFILLER_49_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14813_ _10460_/X _14813_/D VGND VGND VPWR VPWR _14813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14744_ _10721_/X _14744_/D VGND VGND VPWR VPWR _14744_/Q sky130_fd_sc_hd__dfxtp_1
X_11956_ _11976_/A VGND VGND VPWR VPWR _11956_/X sky130_fd_sc_hd__buf_1
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10907_ _10909_/A VGND VGND VPWR VPWR _10907_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11887_ _11896_/A VGND VGND VPWR VPWR _11887_/X sky130_fd_sc_hd__buf_1
X_14675_ _11005_/X _14675_/D VGND VGND VPWR VPWR _14675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater20 _13950_/S1 VGND VGND VPWR VPWR _07541_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_60_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13626_ _13625_/X _14310_/D _15506_/Q VGND VGND VPWR VPWR _13626_/X sky130_fd_sc_hd__mux2_2
X_10838_ _10838_/A _10838_/B VGND VGND VPWR VPWR _10851_/A sky130_fd_sc_hd__or2_2
Xrepeater31 _14399_/Q VGND VGND VPWR VPWR _13945_/S0 sky130_fd_sc_hd__clkbuf_16
Xrepeater42 _14396_/Q VGND VGND VPWR VPWR _14210_/S1 sky130_fd_sc_hd__clkbuf_16
Xrepeater53 _14387_/Q VGND VGND VPWR VPWR _13648_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_9_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10769_ _10769_/A VGND VGND VPWR VPWR _10769_/X sky130_fd_sc_hd__clkbuf_1
X_13557_ _13556_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13557_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12508_ _12492_/A _12507_/A _12951_/B _12507_/Y VGND VGND VPWR VPWR _12513_/A sky130_fd_sc_hd__o22a_1
X_13488_ _13856_/X _13861_/X _13521_/S VGND VGND VPWR VPWR _13488_/X sky130_fd_sc_hd__mux2_1
X_12439_ _15557_/Q VGND VGND VPWR VPWR _12902_/B sky130_fd_sc_hd__buf_1
X_15227_ _08816_/X _15227_/D VGND VGND VPWR VPWR _15227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15158_ _09083_/X _15158_/D VGND VGND VPWR VPWR _15158_/Q sky130_fd_sc_hd__dfxtp_1
X_14109_ _14837_/Q _14869_/Q _14901_/Q _14933_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14109_/X sky130_fd_sc_hd__mux4_2
XFILLER_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15089_ _09361_/X _15089_/D VGND VGND VPWR VPWR _15089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07980_ _07986_/A VGND VGND VPWR VPWR _07980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09650_ _15020_/Q _09641_/X _09649_/X _09645_/X VGND VGND VPWR VPWR _15020_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08601_ _08603_/A VGND VGND VPWR VPWR _08601_/X sky130_fd_sc_hd__clkbuf_1
X_09581_ _15033_/Q _09577_/X _09579_/X _09580_/X VGND VGND VPWR VPWR _15033_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08532_ _08542_/A VGND VGND VPWR VPWR _08532_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08463_ _08463_/A VGND VGND VPWR VPWR _08463_/X sky130_fd_sc_hd__buf_1
XFILLER_50_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07414_ _07415_/A _13575_/X VGND VGND VPWR VPWR _15580_/D sky130_fd_sc_hd__and2_1
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08394_ _14328_/Q VGND VGND VPWR VPWR _10707_/A sky130_fd_sc_hd__buf_1
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07345_ _07353_/A _07345_/B VGND VGND VPWR VPWR _15600_/D sky130_fd_sc_hd__nor2_1
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_30_clk _14397_/CLK VGND VGND VPWR VPWR _15458_/CLK sky130_fd_sc_hd__clkbuf_16
X_07276_ _07278_/A _07276_/B VGND VGND VPWR VPWR _15618_/D sky130_fd_sc_hd__nor2_1
XFILLER_136_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09015_ _09021_/A VGND VGND VPWR VPWR _09015_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09917_ _09917_/A VGND VGND VPWR VPWR _09952_/A sky130_fd_sc_hd__buf_1
XFILLER_59_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09848_ _14969_/Q _09846_/X _09579_/X _09847_/X VGND VGND VPWR VPWR _14969_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09779_ _09798_/A VGND VGND VPWR VPWR _09779_/X sky130_fd_sc_hd__buf_1
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11810_ _11818_/A VGND VGND VPWR VPWR _11810_/X sky130_fd_sc_hd__clkbuf_1
X_12790_ _12775_/X _12788_/X _12789_/X _13285_/X _12710_/X VGND VGND VPWR VPWR _12790_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11741_ _14484_/Q _11733_/X _11498_/X _11735_/X VGND VGND VPWR VPWR _14484_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11672_ _11678_/A VGND VGND VPWR VPWR _11672_/X sky130_fd_sc_hd__clkbuf_1
X_14460_ _11824_/X _14460_/D VGND VGND VPWR VPWR _14460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13411_ _12737_/A _12730_/A _13418_/S VGND VGND VPWR VPWR _13411_/X sky130_fd_sc_hd__mux2_1
X_10623_ _10625_/A VGND VGND VPWR VPWR _10623_/X sky130_fd_sc_hd__clkbuf_1
X_14391_ _14391_/CLK instruction[28] VGND VGND VPWR VPWR _14391_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_21_clk _14328_/CLK VGND VGND VPWR VPWR _15591_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13342_ _13341_/X _13350_/X _13393_/S VGND VGND VPWR VPWR _13342_/X sky130_fd_sc_hd__mux2_1
X_10554_ _14786_/Q _10550_/X _10297_/X _10553_/X VGND VGND VPWR VPWR _14786_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13273_ _13272_/X _12376_/X _15565_/Q VGND VGND VPWR VPWR _13273_/X sky130_fd_sc_hd__mux2_1
X_10485_ _10516_/A VGND VGND VPWR VPWR _10506_/A sky130_fd_sc_hd__buf_2
X_12224_ _15562_/Q VGND VGND VPWR VPWR _12815_/A sky130_fd_sc_hd__inv_2
X_15012_ _09689_/X _15012_/D VGND VGND VPWR VPWR _15012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12155_ _15575_/Q VGND VGND VPWR VPWR _12155_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11106_ _11111_/A VGND VGND VPWR VPWR _11106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12086_ _12086_/A VGND VGND VPWR VPWR _12087_/B sky130_fd_sc_hd__inv_2
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11037_ _11046_/A VGND VGND VPWR VPWR _11037_/X sky130_fd_sc_hd__buf_1
XFILLER_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12988_ _15518_/Q _12575_/A _07633_/B _07387_/A _12987_/X VGND VGND VPWR VPWR _12988_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_18_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14727_ _10811_/X _14727_/D VGND VGND VPWR VPWR _14727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11939_ _11941_/A VGND VGND VPWR VPWR _11939_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14658_ _11060_/X _14658_/D VGND VGND VPWR VPWR _14658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13609_ _13608_/X _07326_/Y _13649_/S VGND VGND VPWR VPWR _13609_/X sky130_fd_sc_hd__mux2_1
X_14589_ _11340_/X _14589_/D VGND VGND VPWR VPWR _14589_/Q sky130_fd_sc_hd__dfxtp_1
X_07130_ _13114_/X VGND VGND VPWR VPWR _07258_/B sky130_fd_sc_hd__inv_2
XFILLER_119_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07963_ _07963_/A VGND VGND VPWR VPWR _07963_/X sky130_fd_sc_hd__clkbuf_2
X_09702_ _09702_/A VGND VGND VPWR VPWR _09702_/X sky130_fd_sc_hd__buf_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07894_ _07889_/A _07889_/B _07893_/X _07889_/Y VGND VGND VPWR VPWR _15433_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09633_ _15023_/Q _09625_/X _09632_/X _09628_/X VGND VGND VPWR VPWR _15023_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09564_ _10328_/A VGND VGND VPWR VPWR _09564_/X sky130_fd_sc_hd__buf_1
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08515_ _14309_/Q VGND VGND VPWR VPWR _10808_/A sky130_fd_sc_hd__buf_1
XFILLER_24_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09495_ _09495_/A VGND VGND VPWR VPWR _09495_/X sky130_fd_sc_hd__clkbuf_1
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08446_ _14320_/Q VGND VGND VPWR VPWR _10750_/A sky130_fd_sc_hd__buf_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08377_ _09176_/A VGND VGND VPWR VPWR _08377_/X sky130_fd_sc_hd__buf_1
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07328_ _07361_/A VGND VGND VPWR VPWR _07337_/A sky130_fd_sc_hd__buf_1
XFILLER_149_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07259_ _07260_/A _07259_/B VGND VGND VPWR VPWR _15629_/D sky130_fd_sc_hd__nor2_1
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10270_ _10270_/A VGND VGND VPWR VPWR _10931_/A sky130_fd_sc_hd__buf_1
XFILLER_118_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13960_ _14948_/Q _15044_/Q _15012_/Q _15076_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13960_/X sky130_fd_sc_hd__mux4_2
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12911_ _12155_/X _12712_/X _12708_/A _12709_/A VGND VGND VPWR VPWR _12914_/B sky130_fd_sc_hd__o22a_1
XFILLER_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13891_ _13887_/X _13888_/X _13889_/X _13890_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13891_/X sky130_fd_sc_hd__mux4_2
X_15630_ _15663_/CLK _15630_/D VGND VGND VPWR VPWR pc[25] sky130_fd_sc_hd__dfxtp_2
XFILLER_64_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12842_ _15534_/Q VGND VGND VPWR VPWR _12842_/X sky130_fd_sc_hd__buf_1
XFILLER_64_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15561_ _15566_/CLK _15561_/D VGND VGND VPWR VPWR _15561_/Q sky130_fd_sc_hd__dfxtp_4
X_12773_ _12773_/A VGND VGND VPWR VPWR _12785_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14512_ _11641_/X _14512_/D VGND VGND VPWR VPWR _14512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11724_ _14489_/Q _11722_/X _11475_/X _11723_/X VGND VGND VPWR VPWR _14489_/D sky130_fd_sc_hd__a22o_1
X_15492_ _15579_/CLK _15492_/D VGND VGND VPWR VPWR wdata[18] sky130_fd_sc_hd__dfxtp_2
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11655_ _14509_/Q _11652_/X _11528_/X _11654_/X VGND VGND VPWR VPWR _14509_/D sky130_fd_sc_hd__a22o_1
X_14443_ _11883_/X _14443_/D VGND VGND VPWR VPWR _14443_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10606_ _10606_/A VGND VGND VPWR VPWR _10606_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14374_ _14385_/CLK instruction[3] VGND VGND VPWR VPWR _14374_/Q sky130_fd_sc_hd__dfxtp_2
X_11586_ _14528_/Q _11578_/X _11443_/X _11581_/X VGND VGND VPWR VPWR _14528_/D sky130_fd_sc_hd__a22o_1
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13325_ _13324_/X _13337_/X _13408_/S VGND VGND VPWR VPWR _13325_/X sky130_fd_sc_hd__mux2_1
X_10537_ _14791_/Q _10535_/X _10419_/X _10536_/X VGND VGND VPWR VPWR _14791_/D sky130_fd_sc_hd__a22o_1
XFILLER_127_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13256_ _13257_/X _12850_/A _13393_/S VGND VGND VPWR VPWR _13256_/X sky130_fd_sc_hd__mux2_2
X_10468_ _10470_/A VGND VGND VPWR VPWR _10468_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12207_ _12275_/A _12275_/B VGND VGND VPWR VPWR _12207_/Y sky130_fd_sc_hd__nor2_1
X_13187_ _12388_/X _12395_/A _13418_/S VGND VGND VPWR VPWR _13187_/X sky130_fd_sc_hd__mux2_1
X_10399_ _10399_/A VGND VGND VPWR VPWR _10399_/X sky130_fd_sc_hd__buf_1
XFILLER_123_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12138_ _12287_/A VGND VGND VPWR VPWR _12138_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_150_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12069_ _12164_/A VGND VGND VPWR VPWR _12092_/A sky130_fd_sc_hd__buf_1
XFILLER_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08300_ _08304_/A VGND VGND VPWR VPWR _08300_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09280_ _15110_/Q _09274_/X _09279_/X _09276_/X VGND VGND VPWR VPWR _15110_/D sky130_fd_sc_hd__a22o_1
X_08231_ _15362_/Q _08227_/X _07929_/X _08230_/X VGND VGND VPWR VPWR _15362_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08162_ _08180_/A VGND VGND VPWR VPWR _08169_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07113_ _07209_/A VGND VGND VPWR VPWR _07291_/A sky130_fd_sc_hd__buf_1
XFILLER_107_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08093_ _08097_/A VGND VGND VPWR VPWR _08093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08995_ _15184_/Q _08993_/X _08865_/X _08994_/X VGND VGND VPWR VPWR _15184_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07946_ _07956_/A VGND VGND VPWR VPWR _07946_/X sky130_fd_sc_hd__clkbuf_1
X_07877_ _07874_/X _07884_/B _07884_/A _07733_/A VGND VGND VPWR VPWR _07878_/B sky130_fd_sc_hd__a31o_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09616_ _10755_/A VGND VGND VPWR VPWR _10371_/A sky130_fd_sc_hd__buf_1
XFILLER_71_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09547_ _09547_/A VGND VGND VPWR VPWR _09644_/A sky130_fd_sc_hd__buf_2
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ _09478_/A VGND VGND VPWR VPWR _09499_/A sky130_fd_sc_hd__buf_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08429_ _08467_/A VGND VGND VPWR VPWR _08429_/X sky130_fd_sc_hd__buf_1
XFILLER_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11440_ _11520_/A VGND VGND VPWR VPWR _11469_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11371_ _11373_/A VGND VGND VPWR VPWR _11371_/X sky130_fd_sc_hd__clkbuf_1
X_13110_ _15656_/Q data_address[21] _15667_/Q VGND VGND VPWR VPWR _13110_/X sky130_fd_sc_hd__mux2_1
X_10322_ _10334_/A VGND VGND VPWR VPWR _10331_/A sky130_fd_sc_hd__buf_1
XFILLER_125_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14090_ _14967_/Q _15063_/Q _15031_/Q _15095_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14090_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13041_ wdata[14] rdata[14] ren VGND VGND VPWR VPWR _14318_/D sky130_fd_sc_hd__mux2_1
X_10253_ _10255_/A VGND VGND VPWR VPWR _10253_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10184_ _10194_/A VGND VGND VPWR VPWR _10197_/A sky130_fd_sc_hd__inv_2
XFILLER_132_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14992_ _09766_/X _14992_/D VGND VGND VPWR VPWR _14992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13943_ _14661_/Q _15237_/Q _14725_/Q _14693_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13943_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13874_ _15180_/Q _15148_/Q _14764_/Q _14796_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13874_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15613_ _15646_/CLK _15613_/D VGND VGND VPWR VPWR pc[8] sky130_fd_sc_hd__dfxtp_2
X_12825_ _12825_/A VGND VGND VPWR VPWR _12825_/X sky130_fd_sc_hd__buf_1
XFILLER_50_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15544_ _15544_/CLK _15544_/D VGND VGND VPWR VPWR _15544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12756_ _12758_/A _12758_/B _12727_/X VGND VGND VPWR VPWR _12756_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11707_ _11716_/A VGND VGND VPWR VPWR _11712_/A sky130_fd_sc_hd__buf_1
X_15475_ _15521_/CLK _15475_/D VGND VGND VPWR VPWR wdata[1] sky130_fd_sc_hd__dfxtp_2
X_12687_ _12686_/X _12209_/X _12279_/X VGND VGND VPWR VPWR _12735_/B sky130_fd_sc_hd__o21ai_1
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14426_ _11941_/X _14426_/D VGND VGND VPWR VPWR _14426_/Q sky130_fd_sc_hd__dfxtp_1
X_11638_ _11638_/A VGND VGND VPWR VPWR _11638_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14357_ _15654_/CLK pc[18] VGND VGND VPWR VPWR _14357_/Q sky130_fd_sc_hd__dfxtp_1
X_11569_ _11569_/A VGND VGND VPWR VPWR _11569_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13308_ _13307_/X _13312_/X _13393_/S VGND VGND VPWR VPWR _13308_/X sky130_fd_sc_hd__mux2_1
X_14288_ _14499_/Q _14467_/Q _14435_/Q _14403_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14288_/X sky130_fd_sc_hd__mux4_1
X_13239_ _13240_/X _13264_/X _15563_/Q VGND VGND VPWR VPWR _13239_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07800_ _07800_/A VGND VGND VPWR VPWR _07800_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08780_ _09700_/A _11576_/A VGND VGND VPWR VPWR _08796_/A sky130_fd_sc_hd__or2_2
XFILLER_38_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07731_ _07731_/A VGND VGND VPWR VPWR _07731_/X sky130_fd_sc_hd__buf_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07662_ _07658_/A _13122_/X _07660_/X _07661_/Y VGND VGND VPWR VPWR _07789_/A sky130_fd_sc_hd__o22a_1
XFILLER_92_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09401_ _15077_/Q _09395_/X _09284_/X _09396_/X VGND VGND VPWR VPWR _15077_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07593_ _07595_/A _13073_/X VGND VGND VPWR VPWR _15488_/D sky130_fd_sc_hd__and2_1
XFILLER_80_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09332_ _15098_/Q _09326_/X _09192_/X _09327_/X VGND VGND VPWR VPWR _15098_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09263_ _09263_/A VGND VGND VPWR VPWR _09263_/X sky130_fd_sc_hd__buf_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08214_ _08216_/A VGND VGND VPWR VPWR _08214_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09194_ _09199_/A VGND VGND VPWR VPWR _09194_/X sky130_fd_sc_hd__clkbuf_1
X_08145_ _15385_/Q _08143_/X _07983_/X _08144_/X VGND VGND VPWR VPWR _15385_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08076_ _08082_/A VGND VGND VPWR VPWR _08076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08978_ _08980_/A VGND VGND VPWR VPWR _08978_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07929_ _07929_/A VGND VGND VPWR VPWR _07929_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10940_ _14694_/Q _10936_/X _10819_/X _10937_/X VGND VGND VPWR VPWR _14694_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10871_ _10901_/A VGND VGND VPWR VPWR _10892_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12610_ _12610_/A VGND VGND VPWR VPWR _12610_/X sky130_fd_sc_hd__buf_4
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ _13589_/X _14319_/D _15506_/Q VGND VGND VPWR VPWR _13590_/X sky130_fd_sc_hd__mux2_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12541_ _15464_/Q _12541_/B VGND VGND VPWR VPWR wen sky130_fd_sc_hd__and2_2
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15260_ _08692_/X _15260_/D VGND VGND VPWR VPWR _15260_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12472_ _12616_/A VGND VGND VPWR VPWR _12472_/X sky130_fd_sc_hd__clkbuf_2
X_14211_ _14207_/X _14208_/X _14209_/X _14210_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14211_/X sky130_fd_sc_hd__mux4_2
X_11423_ _14564_/Q _11319_/A _11198_/X _11322_/A VGND VGND VPWR VPWR _14564_/D sky130_fd_sc_hd__a22o_1
X_15191_ _08968_/X _15191_/D VGND VGND VPWR VPWR _15191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ _15217_/Q _14545_/Q _14993_/Q _15409_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14142_/X sky130_fd_sc_hd__mux4_1
X_11354_ _11354_/A VGND VGND VPWR VPWR _11354_/X sky130_fd_sc_hd__buf_1
XFILLER_137_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10305_ _10346_/A VGND VGND VPWR VPWR _10334_/A sky130_fd_sc_hd__clkbuf_2
X_14073_ _14680_/Q _15256_/Q _14744_/Q _14712_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14073_/X sky130_fd_sc_hd__mux4_2
XFILLER_4_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11285_ _11285_/A VGND VGND VPWR VPWR _11304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10236_ _10236_/A VGND VGND VPWR VPWR _10236_/X sky130_fd_sc_hd__clkbuf_1
X_13024_ _14368_/Q VGND VGND VPWR VPWR _13024_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10167_ _10167_/A VGND VGND VPWR VPWR _10167_/X sky130_fd_sc_hd__buf_1
XFILLER_86_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14975_ _09822_/X _14975_/D VGND VGND VPWR VPWR _14975_/Q sky130_fd_sc_hd__dfxtp_1
X_10098_ _10107_/A VGND VGND VPWR VPWR _10098_/X sky130_fd_sc_hd__buf_1
X_13926_ _13922_/X _13923_/X _13924_/X _13925_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13926_/X sky130_fd_sc_hd__mux4_2
XFILLER_75_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13857_ _14638_/Q _14606_/Q _14574_/Q _15374_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13857_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12808_ _12812_/A _12812_/B _12328_/X VGND VGND VPWR VPWR _12808_/X sky130_fd_sc_hd__o21a_1
X_13788_ _14517_/Q _14485_/Q _14453_/Q _14421_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13788_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15527_ _15527_/CLK _15527_/D VGND VGND VPWR VPWR _15527_/Q sky130_fd_sc_hd__dfxtp_1
X_12739_ _12739_/A VGND VGND VPWR VPWR _12879_/A sky130_fd_sc_hd__inv_2
XFILLER_148_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15458_ _15458_/CLK _15458_/D VGND VGND VPWR VPWR data_address[31] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14409_ _11999_/X _14409_/D VGND VGND VPWR VPWR _14409_/Q sky130_fd_sc_hd__dfxtp_1
X_15389_ _08129_/X _15389_/D VGND VGND VPWR VPWR _15389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09950_ _10320_/A VGND VGND VPWR VPWR _09950_/X sky130_fd_sc_hd__buf_1
XFILLER_98_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08901_ _09271_/A VGND VGND VPWR VPWR _08901_/X sky130_fd_sc_hd__buf_1
X_09881_ _09885_/A VGND VGND VPWR VPWR _09881_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08832_ _08846_/A VGND VGND VPWR VPWR _08843_/A sky130_fd_sc_hd__buf_2
XFILLER_98_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08763_ _08763_/A VGND VGND VPWR VPWR _08763_/X sky130_fd_sc_hd__buf_1
XFILLER_85_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07714_ _07647_/A _13137_/X _07647_/A _13137_/X VGND VGND VPWR VPWR _07861_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08694_ _08703_/A VGND VGND VPWR VPWR _08694_/X sky130_fd_sc_hd__buf_1
XFILLER_26_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07645_ _07715_/A VGND VGND VPWR VPWR _07679_/A sky130_fd_sc_hd__buf_1
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07576_ _07577_/A _13084_/X VGND VGND VPWR VPWR _15499_/D sky130_fd_sc_hd__and2_1
X_09315_ _15103_/Q _09311_/X _09170_/X _09314_/X VGND VGND VPWR VPWR _15103_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09246_ _15118_/Q _09235_/X _09245_/X _09237_/X VGND VGND VPWR VPWR _15118_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09177_ _15134_/Q _09169_/X _09176_/X _09173_/X VGND VGND VPWR VPWR _15134_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08128_ _15390_/Q _08122_/X _07958_/X _08125_/X VGND VGND VPWR VPWR _15390_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08059_ _08059_/A VGND VGND VPWR VPWR _08059_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11070_ _11070_/A VGND VGND VPWR VPWR _11070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10021_ _14926_/Q _10011_/X _10020_/X _10013_/X VGND VGND VPWR VPWR _14926_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14760_ _10643_/X _14760_/D VGND VGND VPWR VPWR _14760_/Q sky130_fd_sc_hd__dfxtp_1
X_11972_ _14417_/Q _11966_/X _08026_/A _11967_/X VGND VGND VPWR VPWR _14417_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13711_ _13707_/X _13708_/X _13709_/X _13710_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13711_/X sky130_fd_sc_hd__mux4_1
X_10923_ _10929_/A VGND VGND VPWR VPWR _10923_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14691_ _10946_/X _14691_/D VGND VGND VPWR VPWR _14691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13642_ _13641_/X _14306_/D _15506_/Q VGND VGND VPWR VPWR _13642_/X sky130_fd_sc_hd__mux2_1
X_10854_ _10854_/A VGND VGND VPWR VPWR _10915_/A sky130_fd_sc_hd__buf_4
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _13572_/X _13581_/A1 _13641_/S VGND VGND VPWR VPWR _13573_/X sky130_fd_sc_hd__mux2_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10785_ _14733_/Q _10780_/X _10782_/X _10784_/X VGND VGND VPWR VPWR _14733_/D sky130_fd_sc_hd__a22o_1
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15312_ _08462_/X _15312_/D VGND VGND VPWR VPWR _15312_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12524_ _12524_/A VGND VGND VPWR VPWR _12962_/A sky130_fd_sc_hd__buf_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15243_ _08750_/X _15243_/D VGND VGND VPWR VPWR _15243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12455_ _12428_/X _12442_/X _12443_/Y _12454_/Y VGND VGND VPWR VPWR _12455_/X sky130_fd_sc_hd__a31o_1
X_11406_ _14570_/Q _11404_/X _11174_/X _11405_/X VGND VGND VPWR VPWR _14570_/D sky130_fd_sc_hd__a22o_1
X_15174_ _09028_/X _15174_/D VGND VGND VPWR VPWR _15174_/Q sky130_fd_sc_hd__dfxtp_1
X_12386_ _15587_/Q VGND VGND VPWR VPWR _12386_/Y sky130_fd_sc_hd__inv_2
X_14125_ _15123_/Q _15347_/Q _15315_/Q _15283_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14125_/X sky130_fd_sc_hd__mux4_1
X_11337_ _11337_/A VGND VGND VPWR VPWR _11342_/A sky130_fd_sc_hd__buf_1
XFILLER_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14056_ _14052_/X _14053_/X _14054_/X _14055_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14056_/X sky130_fd_sc_hd__mux4_2
X_11268_ _14610_/Q _11264_/X _11138_/X _11265_/X VGND VGND VPWR VPWR _14610_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13007_ _14351_/Q VGND VGND VPWR VPWR _13007_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10219_ _14873_/Q _10217_/X _09973_/X _10218_/X VGND VGND VPWR VPWR _14873_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11199_ _14628_/Q _11064_/A _11198_/X _11068_/A VGND VGND VPWR VPWR _14628_/D sky130_fd_sc_hd__a22o_1
XFILLER_121_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14958_ _09883_/X _14958_/D VGND VGND VPWR VPWR _14958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13909_ _14825_/Q _14857_/Q _14889_/Q _14921_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13909_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14889_ _10160_/X _14889_/D VGND VGND VPWR VPWR _14889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07430_ _07432_/A _13619_/X VGND VGND VPWR VPWR _15569_/D sky130_fd_sc_hd__and2_1
XFILLER_63_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07361_ _07361_/A VGND VGND VPWR VPWR _07377_/A sky130_fd_sc_hd__buf_1
X_09100_ _09120_/A VGND VGND VPWR VPWR _09105_/A sky130_fd_sc_hd__buf_1
XFILLER_31_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07292_ _14394_/Q VGND VGND VPWR VPWR _07313_/B sky130_fd_sc_hd__inv_2
X_09031_ _15173_/Q _09025_/X _08913_/X _09026_/X VGND VGND VPWR VPWR _15173_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09933_ _09933_/A VGND VGND VPWR VPWR _09933_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09864_ _14965_/Q _09856_/X _09601_/X _09858_/X VGND VGND VPWR VPWR _14965_/D sky130_fd_sc_hd__a22o_1
XFILLER_98_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08815_ _15228_/Q _08812_/X _08813_/X _08814_/X VGND VGND VPWR VPWR _15228_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09795_ _09817_/A VGND VGND VPWR VPWR _09802_/A sky130_fd_sc_hd__buf_1
X_08746_ _08746_/A VGND VGND VPWR VPWR _08765_/A sky130_fd_sc_hd__buf_1
XFILLER_38_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_207 _13506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_218 _11190_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_229 _08743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08677_ _08677_/A VGND VGND VPWR VPWR _08741_/A sky130_fd_sc_hd__buf_4
XFILLER_54_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07628_ _07630_/A _07628_/B VGND VGND VPWR VPWR _15470_/D sky130_fd_sc_hd__nor2_1
X_07559_ _07559_/A _07559_/B _07559_/C _07559_/D VGND VGND VPWR VPWR _07559_/X sky130_fd_sc_hd__or4_4
XFILLER_41_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10570_ _10574_/A VGND VGND VPWR VPWR _10570_/X sky130_fd_sc_hd__clkbuf_1
X_09229_ _15122_/Q _09223_/X _09228_/X _09225_/X VGND VGND VPWR VPWR _15122_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12240_ _12806_/A _12238_/A _12239_/X VGND VGND VPWR VPWR _12264_/A sky130_fd_sc_hd__o21a_1
XFILLER_147_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12171_ _12271_/A VGND VGND VPWR VPWR _12725_/A sky130_fd_sc_hd__buf_1
XFILLER_123_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11122_ _11162_/A VGND VGND VPWR VPWR _11149_/A sky130_fd_sc_hd__buf_2
XFILLER_122_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11053_ _14661_/Q _11046_/X _10824_/X _11047_/X VGND VGND VPWR VPWR _14661_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10004_ _14930_/Q _09998_/X _10003_/X _10000_/X VGND VGND VPWR VPWR _14930_/D sky130_fd_sc_hd__a22o_1
XFILLER_131_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14812_ _10464_/X _14812_/D VGND VGND VPWR VPWR _14812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14743_ _10726_/X _14743_/D VGND VGND VPWR VPWR _14743_/Q sky130_fd_sc_hd__dfxtp_1
X_11955_ _11985_/A VGND VGND VPWR VPWR _11976_/A sky130_fd_sc_hd__buf_2
XFILLER_45_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10906_ _14704_/Q _10904_/X _10766_/X _10905_/X VGND VGND VPWR VPWR _14704_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14674_ _11010_/X _14674_/D VGND VGND VPWR VPWR _14674_/Q sky130_fd_sc_hd__dfxtp_1
X_11886_ _11895_/A VGND VGND VPWR VPWR _11886_/X sky130_fd_sc_hd__buf_1
Xrepeater10 _15562_/Q VGND VGND VPWR VPWR _13415_/S sky130_fd_sc_hd__clkbuf_16
X_13625_ _13624_/X _07348_/Y _13641_/S VGND VGND VPWR VPWR _13625_/X sky130_fd_sc_hd__mux2_1
X_10837_ _10847_/A VGND VGND VPWR VPWR _10837_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater21 _14400_/Q VGND VGND VPWR VPWR _13950_/S1 sky130_fd_sc_hd__clkbuf_16
XFILLER_20_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater32 _14266_/S1 VGND VGND VPWR VPWR _14286_/S1 sky130_fd_sc_hd__clkbuf_16
Xrepeater43 _14055_/S0 VGND VGND VPWR VPWR _14283_/S0 sky130_fd_sc_hd__clkbuf_16
Xrepeater54 _14386_/Q VGND VGND VPWR VPWR _13521_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_13_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13556_ _14056_/X _14061_/X _14387_/Q VGND VGND VPWR VPWR _13556_/X sky130_fd_sc_hd__mux2_2
X_10768_ _14736_/Q _10764_/X _10766_/X _10767_/X VGND VGND VPWR VPWR _14736_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12507_ _12507_/A VGND VGND VPWR VPWR _12507_/Y sky130_fd_sc_hd__inv_2
X_13487_ _13486_/X _13071_/X _14336_/Q VGND VGND VPWR VPWR _13487_/X sky130_fd_sc_hd__mux2_1
X_10699_ _14749_/Q _10682_/X _10698_/X _10687_/X VGND VGND VPWR VPWR _14749_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15226_ _08821_/X _15226_/D VGND VGND VPWR VPWR _15226_/Q sky130_fd_sc_hd__dfxtp_1
X_12438_ _15589_/Q _12347_/A _12902_/A _12505_/A VGND VGND VPWR VPWR _12440_/A sky130_fd_sc_hd__o22a_1
XFILLER_114_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15157_ _09090_/X _15157_/D VGND VGND VPWR VPWR _15157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12369_ _12369_/A VGND VGND VPWR VPWR _12670_/A sky130_fd_sc_hd__buf_1
XFILLER_113_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14108_ _14517_/Q _14485_/Q _14453_/Q _14421_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14108_/X sky130_fd_sc_hd__mux4_1
X_15088_ _09364_/X _15088_/D VGND VGND VPWR VPWR _15088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14039_ _14844_/Q _14876_/Q _14908_/Q _14940_/Q _14395_/Q _14060_/S1 VGND VGND VPWR
+ VPWR _14039_/X sky130_fd_sc_hd__mux4_2
XFILLER_68_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08600_ _15286_/Q _08597_/X _08427_/X _08599_/X VGND VGND VPWR VPWR _15286_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09580_ _09580_/A VGND VGND VPWR VPWR _09580_/X sky130_fd_sc_hd__buf_1
X_08531_ _08531_/A VGND VGND VPWR VPWR _08542_/A sky130_fd_sc_hd__buf_2
XFILLER_36_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08462_ _08469_/A VGND VGND VPWR VPWR _08462_/X sky130_fd_sc_hd__clkbuf_1
X_07413_ _07415_/A _13571_/X VGND VGND VPWR VPWR _15581_/D sky130_fd_sc_hd__and2_1
X_08393_ _08393_/A VGND VGND VPWR VPWR _08393_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07344_ _07361_/A VGND VGND VPWR VPWR _07353_/A sky130_fd_sc_hd__buf_1
XFILLER_148_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07275_ _07283_/A VGND VGND VPWR VPWR _07278_/A sky130_fd_sc_hd__buf_1
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09014_ _09023_/A VGND VGND VPWR VPWR _09021_/A sky130_fd_sc_hd__buf_1
XFILLER_145_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09916_ _14948_/Q _09812_/A _09691_/X _09815_/A VGND VGND VPWR VPWR _14948_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09847_ _09847_/A VGND VGND VPWR VPWR _09847_/X sky130_fd_sc_hd__buf_1
XFILLER_74_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09778_ _09778_/A VGND VGND VPWR VPWR _09798_/A sky130_fd_sc_hd__buf_1
XFILLER_27_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08729_ _08731_/A VGND VGND VPWR VPWR _08729_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11740_ _11742_/A VGND VGND VPWR VPWR _11740_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11671_ _11680_/A VGND VGND VPWR VPWR _11678_/A sky130_fd_sc_hd__buf_1
XFILLER_53_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13410_ _12709_/X _12703_/A _13418_/S VGND VGND VPWR VPWR _13410_/X sky130_fd_sc_hd__mux2_1
X_10622_ _14767_/Q _10616_/X _10383_/X _10617_/X VGND VGND VPWR VPWR _14767_/D sky130_fd_sc_hd__a22o_1
X_14390_ _15648_/CLK instruction[27] VGND VGND VPWR VPWR _14390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13341_ _13340_/X _13353_/X _13408_/S VGND VGND VPWR VPWR _13341_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10553_ _10553_/A VGND VGND VPWR VPWR _10553_/X sky130_fd_sc_hd__buf_1
XFILLER_10_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13272_ _13350_/X _13347_/X _13393_/S VGND VGND VPWR VPWR _13272_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10484_ _10505_/A VGND VGND VPWR VPWR _10484_/X sky130_fd_sc_hd__buf_1
XFILLER_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15011_ _09693_/X _15011_/D VGND VGND VPWR VPWR _15011_/Q sky130_fd_sc_hd__dfxtp_1
X_12223_ _12223_/A VGND VGND VPWR VPWR _12885_/A sky130_fd_sc_hd__buf_1
XFILLER_135_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12154_ _12160_/A VGND VGND VPWR VPWR _12709_/A sky130_fd_sc_hd__buf_1
X_11105_ _14650_/Q _11094_/X _11104_/X _11096_/X VGND VGND VPWR VPWR _14650_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12085_ _12079_/X _12082_/X _12591_/A _12084_/X VGND VGND VPWR VPWR _12086_/A sky130_fd_sc_hd__o22a_1
XFILLER_1_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11036_ _11036_/A VGND VGND VPWR VPWR _11036_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12987_ _07630_/B _14397_/Q _15516_/Q _12572_/A VGND VGND VPWR VPWR _12987_/X sky130_fd_sc_hd__o22a_1
XFILLER_33_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14726_ _10817_/X _14726_/D VGND VGND VPWR VPWR _14726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11938_ _14428_/Q _11936_/X _07968_/A _11937_/X VGND VGND VPWR VPWR _14428_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14657_ _11070_/X _14657_/D VGND VGND VPWR VPWR _14657_/Q sky130_fd_sc_hd__dfxtp_1
X_11869_ _14447_/Q _11865_/X _08036_/A _11866_/X VGND VGND VPWR VPWR _14447_/D sky130_fd_sc_hd__a22o_1
X_13608_ _14186_/X _14191_/X _13648_/S VGND VGND VPWR VPWR _13608_/X sky130_fd_sc_hd__mux2_4
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14588_ _11342_/X _14588_/D VGND VGND VPWR VPWR _14588_/Q sky130_fd_sc_hd__dfxtp_1
X_13539_ _13538_/X _13087_/X _14337_/Q VGND VGND VPWR VPWR _13539_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15209_ _08894_/X _15209_/D VGND VGND VPWR VPWR _15209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07962_ _14330_/Q VGND VGND VPWR VPWR _07963_/A sky130_fd_sc_hd__buf_1
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09701_ _09713_/A VGND VGND VPWR VPWR _09702_/A sky130_fd_sc_hd__buf_1
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07893_ _07893_/A VGND VGND VPWR VPWR _07893_/X sky130_fd_sc_hd__buf_1
XFILLER_56_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09632_ _10383_/A VGND VGND VPWR VPWR _09632_/X sky130_fd_sc_hd__buf_1
XFILLER_55_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09563_ _10702_/A VGND VGND VPWR VPWR _10328_/A sky130_fd_sc_hd__buf_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08514_ _08526_/A VGND VGND VPWR VPWR _08514_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09494_ _15051_/Q _09486_/X _09259_/X _09488_/X VGND VGND VPWR VPWR _15051_/D sky130_fd_sc_hd__a22o_1
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08445_ _08463_/A VGND VGND VPWR VPWR _08445_/X sky130_fd_sc_hd__buf_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08376_ _10690_/A VGND VGND VPWR VPWR _09176_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07327_ _07383_/A VGND VGND VPWR VPWR _07361_/A sky130_fd_sc_hd__buf_1
XFILLER_109_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07258_ _07260_/A _07258_/B VGND VGND VPWR VPWR _15630_/D sky130_fd_sc_hd__nor2_1
XFILLER_125_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07189_ _07251_/B _07179_/B _07188_/X _07180_/Y VGND VGND VPWR VPWR _15665_/D sky130_fd_sc_hd__a211oi_2
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12910_ _12692_/X _12146_/X _12693_/A _12694_/A VGND VGND VPWR VPWR _12941_/A sky130_fd_sc_hd__o22a_1
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13890_ _14955_/Q _15051_/Q _15019_/Q _15083_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13890_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12841_ _12798_/X _12840_/X _12798_/X _12840_/X VGND VGND VPWR VPWR _12841_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_62_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15560_ _15579_/CLK _15560_/D VGND VGND VPWR VPWR _15560_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12772_ _12929_/A _13338_/X VGND VGND VPWR VPWR _12878_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14511_ _11645_/X _14511_/D VGND VGND VPWR VPWR _14511_/Q sky130_fd_sc_hd__dfxtp_1
X_11723_ _11723_/A VGND VGND VPWR VPWR _11723_/X sky130_fd_sc_hd__buf_1
X_15491_ _15597_/CLK _15491_/D VGND VGND VPWR VPWR wdata[17] sky130_fd_sc_hd__dfxtp_2
XFILLER_42_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _11885_/X _14442_/D VGND VGND VPWR VPWR _14442_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11674_/A VGND VGND VPWR VPWR _11654_/X sky130_fd_sc_hd__buf_1
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10605_ _14772_/Q _10597_/X _10363_/X _10599_/X VGND VGND VPWR VPWR _14772_/D sky130_fd_sc_hd__a22o_1
X_14373_ _14381_/CLK instruction[2] VGND VGND VPWR VPWR _14373_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11585_ _11585_/A VGND VGND VPWR VPWR _11585_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13324_ _13385_/X _13384_/X _13415_/S VGND VGND VPWR VPWR _13324_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10536_ _10536_/A VGND VGND VPWR VPWR _10536_/X sky130_fd_sc_hd__buf_1
XFILLER_109_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13255_ _13254_/X _12459_/X _15565_/Q VGND VGND VPWR VPWR _13255_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10467_ _14812_/Q _10465_/X _10328_/X _10466_/X VGND VGND VPWR VPWR _14812_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12206_ _12204_/X _12157_/X _12779_/A _12148_/X VGND VGND VPWR VPWR _12275_/B sky130_fd_sc_hd__o22a_1
XFILLER_89_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13186_ _13187_/X _13197_/X _13415_/S VGND VGND VPWR VPWR _13186_/X sky130_fd_sc_hd__mux2_1
X_10398_ _10398_/A VGND VGND VPWR VPWR _10398_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12137_ _12142_/A VGND VGND VPWR VPWR _12287_/A sky130_fd_sc_hd__buf_1
XFILLER_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12068_ _12156_/A VGND VGND VPWR VPWR _12164_/A sky130_fd_sc_hd__buf_1
XFILLER_38_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11019_ _11023_/A VGND VGND VPWR VPWR _11019_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14709_ _10888_/X _14709_/D VGND VGND VPWR VPWR _14709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08230_ _08230_/A VGND VGND VPWR VPWR _08230_/X sky130_fd_sc_hd__buf_1
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08161_ _08161_/A VGND VGND VPWR VPWR _08180_/A sky130_fd_sc_hd__buf_4
X_07112_ _07182_/A VGND VGND VPWR VPWR _07209_/A sky130_fd_sc_hd__clkbuf_2
X_08092_ _15397_/Q _08077_/X _08091_/X _08080_/X VGND VGND VPWR VPWR _15397_/D sky130_fd_sc_hd__a22o_1
XFILLER_146_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08994_ _08994_/A VGND VGND VPWR VPWR _08994_/X sky130_fd_sc_hd__buf_1
XFILLER_88_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07945_ _15424_/Q _07927_/X _07944_/X _07932_/X VGND VGND VPWR VPWR _15424_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07876_ _07876_/A VGND VGND VPWR VPWR _07884_/A sky130_fd_sc_hd__buf_1
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09615_ _09615_/A VGND VGND VPWR VPWR _09615_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09546_ _10314_/A VGND VGND VPWR VPWR _09546_/X sky130_fd_sc_hd__buf_1
XFILLER_24_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ _15056_/Q _09475_/X _09236_/X _09476_/X VGND VGND VPWR VPWR _15056_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08428_ _08486_/A VGND VGND VPWR VPWR _08467_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08359_ _14333_/Q VGND VGND VPWR VPWR _10676_/A sky130_fd_sc_hd__buf_1
XFILLER_137_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11370_ _14581_/Q _11364_/X _11126_/X _11366_/X VGND VGND VPWR VPWR _14581_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10321_ _14846_/Q _10313_/X _10320_/X _10317_/X VGND VGND VPWR VPWR _14846_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13040_ wdata[13] rdata[13] ren VGND VGND VPWR VPWR _14317_/D sky130_fd_sc_hd__mux2_1
X_10252_ _14863_/Q _10247_/X _10016_/X _10248_/X VGND VGND VPWR VPWR _14863_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10183_ _10183_/A VGND VGND VPWR VPWR _10183_/X sky130_fd_sc_hd__buf_1
XFILLER_59_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14991_ _09770_/X _14991_/D VGND VGND VPWR VPWR _14991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13942_ _15205_/Q _14533_/Q _14981_/Q _15397_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13942_/X sky130_fd_sc_hd__mux4_2
XFILLER_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13873_ _14668_/Q _15244_/Q _14732_/Q _14700_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13873_/X sky130_fd_sc_hd__mux4_2
X_15612_ _15648_/CLK _15612_/D VGND VGND VPWR VPWR pc[7] sky130_fd_sc_hd__dfxtp_4
XFILLER_34_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12824_ _12824_/A VGND VGND VPWR VPWR _12824_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15543_ _15544_/CLK _15543_/D VGND VGND VPWR VPWR _15543_/Q sky130_fd_sc_hd__dfxtp_1
X_12755_ _12755_/A VGND VGND VPWR VPWR _12758_/B sky130_fd_sc_hd__buf_1
X_11706_ _14495_/Q _11702_/X _11449_/X _11705_/X VGND VGND VPWR VPWR _14495_/D sky130_fd_sc_hd__a22o_1
X_15474_ _15579_/CLK _15474_/D VGND VGND VPWR VPWR wdata[0] sky130_fd_sc_hd__dfxtp_2
X_12686_ _12747_/A VGND VGND VPWR VPWR _12686_/X sky130_fd_sc_hd__buf_1
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _11945_/X _14425_/D VGND VGND VPWR VPWR _14425_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ _14514_/Q _11633_/X _11506_/X _11634_/X VGND VGND VPWR VPWR _14514_/D sky130_fd_sc_hd__a22o_1
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _15652_/CLK pc[17] VGND VGND VPWR VPWR _14356_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11568_ _14532_/Q _11430_/A _11567_/X _11434_/A VGND VGND VPWR VPWR _14532_/D sky130_fd_sc_hd__a22o_1
X_13307_ _13382_/X _13379_/X _13408_/S VGND VGND VPWR VPWR _13307_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10519_ _10521_/A VGND VGND VPWR VPWR _10519_/X sky130_fd_sc_hd__clkbuf_1
X_14287_ _14627_/Q _14595_/Q _14563_/Q _15363_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14287_/X sky130_fd_sc_hd__mux4_1
X_11499_ _14548_/Q _11488_/X _11498_/X _11491_/X VGND VGND VPWR VPWR _14548_/D sky130_fd_sc_hd__a22o_1
X_13238_ _13239_/X _13286_/X _13393_/S VGND VGND VPWR VPWR _13238_/X sky130_fd_sc_hd__mux2_2
XFILLER_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13169_ _13168_/X _13191_/X _13408_/S VGND VGND VPWR VPWR _13169_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07730_ _13144_/X _07730_/B VGND VGND VPWR VPWR _07731_/A sky130_fd_sc_hd__nor2_1
XFILLER_84_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07661_ _13122_/X VGND VGND VPWR VPWR _07661_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09400_ _09400_/A VGND VGND VPWR VPWR _09400_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07592_ _07596_/A VGND VGND VPWR VPWR _07595_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09331_ _09331_/A VGND VGND VPWR VPWR _09331_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09262_ _09274_/A VGND VGND VPWR VPWR _09262_/X sky130_fd_sc_hd__buf_1
X_08213_ _15364_/Q _08109_/A _08095_/X _08112_/A VGND VGND VPWR VPWR _15364_/D sky130_fd_sc_hd__a22o_1
X_09193_ _15130_/Q _09183_/X _09192_/X _09185_/X VGND VGND VPWR VPWR _15130_/D sky130_fd_sc_hd__a22o_1
X_08144_ _08144_/A VGND VGND VPWR VPWR _08144_/X sky130_fd_sc_hd__buf_1
XFILLER_146_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08075_ _15400_/Q _08062_/X _08074_/X _08065_/X VGND VGND VPWR VPWR _15400_/D sky130_fd_sc_hd__a22o_1
XFILLER_146_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08977_ _15190_/Q _08974_/X _08839_/X _08976_/X VGND VGND VPWR VPWR _15190_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07928_ _14335_/Q VGND VGND VPWR VPWR _07929_/A sky130_fd_sc_hd__buf_1
XFILLER_29_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07859_ _07848_/X _07711_/X _07864_/B VGND VGND VPWR VPWR _07860_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10870_ _14714_/Q _10864_/X _10713_/X _10865_/X VGND VGND VPWR VPWR _14714_/D sky130_fd_sc_hd__a22o_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09529_ _09547_/A VGND VGND VPWR VPWR _09530_/A sky130_fd_sc_hd__buf_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12540_ _15464_/Q _12541_/B VGND VGND VPWR VPWR ren sky130_fd_sc_hd__nor2b_4
XFILLER_24_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12471_ _12500_/A VGND VGND VPWR VPWR _12616_/A sky130_fd_sc_hd__buf_1
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14210_ _14955_/Q _15051_/Q _15019_/Q _15083_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14210_/X sky130_fd_sc_hd__mux4_2
X_11422_ _11422_/A VGND VGND VPWR VPWR _11422_/X sky130_fd_sc_hd__buf_1
X_15190_ _08972_/X _15190_/D VGND VGND VPWR VPWR _15190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14141_ _14137_/X _14138_/X _14139_/X _14140_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14141_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11353_ _11353_/A VGND VGND VPWR VPWR _11353_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10304_ _14849_/Q _10296_/X _10303_/X _10300_/X VGND VGND VPWR VPWR _14849_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14072_ _15224_/Q _14552_/Q _15000_/Q _15416_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14072_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11284_ _11303_/A VGND VGND VPWR VPWR _11284_/X sky130_fd_sc_hd__buf_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13023_ _14367_/Q VGND VGND VPWR VPWR _13023_/Y sky130_fd_sc_hd__inv_2
X_10235_ _14868_/Q _10227_/X _09995_/X _10229_/X VGND VGND VPWR VPWR _14868_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10166_ _10166_/A VGND VGND VPWR VPWR _10166_/X sky130_fd_sc_hd__buf_1
XFILLER_79_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14974_ _09832_/X _14974_/D VGND VGND VPWR VPWR _14974_/Q sky130_fd_sc_hd__dfxtp_1
X_10097_ _10106_/A VGND VGND VPWR VPWR _10097_/X sky130_fd_sc_hd__buf_1
XFILLER_35_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13925_ _15111_/Q _15335_/Q _15303_/Q _15271_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13925_/X sky130_fd_sc_hd__mux4_1
X_13856_ _13852_/X _13853_/X _13854_/X _13855_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13856_/X sky130_fd_sc_hd__mux4_2
X_12807_ _12807_/A VGND VGND VPWR VPWR _12812_/B sky130_fd_sc_hd__buf_1
XFILLER_50_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13787_ _14645_/Q _14613_/Q _14581_/Q _15381_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13787_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10999_ _10999_/A VGND VGND VPWR VPWR _11018_/A sky130_fd_sc_hd__clkbuf_2
X_12738_ _12593_/A _12913_/B _12448_/X VGND VGND VPWR VPWR _12738_/X sky130_fd_sc_hd__o21a_1
X_15526_ _15527_/CLK _15526_/D VGND VGND VPWR VPWR _15526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15457_ _15666_/CLK _15457_/D VGND VGND VPWR VPWR data_address[30] sky130_fd_sc_hd__dfxtp_1
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ _12138_/X _12668_/X _12450_/X _13229_/X _12383_/X VGND VGND VPWR VPWR _12669_/X
+ sky130_fd_sc_hd__o32a_1
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14408_ _12001_/X _14408_/D VGND VGND VPWR VPWR _14408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15388_ _08133_/X _15388_/D VGND VGND VPWR VPWR _15388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14339_ _15601_/CLK pc[0] VGND VGND VPWR VPWR _14339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08900_ _08908_/A VGND VGND VPWR VPWR _08900_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09880_ _09880_/A VGND VGND VPWR VPWR _09885_/A sky130_fd_sc_hd__buf_2
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08831_ _15224_/Q _08825_/X _08830_/X _08827_/X VGND VGND VPWR VPWR _15224_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_opt_7_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR clkbuf_opt_7_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_98_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08762_ _08762_/A VGND VGND VPWR VPWR _08762_/X sky130_fd_sc_hd__buf_1
XFILLER_85_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07713_ _07680_/A _07711_/X _07680_/A _13138_/X VGND VGND VPWR VPWR _07863_/A sky130_fd_sc_hd__a2bb2o_1
X_08693_ _08702_/A VGND VGND VPWR VPWR _08693_/X sky130_fd_sc_hd__buf_1
XFILLER_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07644_ _07660_/A VGND VGND VPWR VPWR _07715_/A sky130_fd_sc_hd__inv_2
XFILLER_26_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07575_ _07577_/A _13085_/X VGND VGND VPWR VPWR _15500_/D sky130_fd_sc_hd__and2_1
XFILLER_53_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09314_ _09336_/A VGND VGND VPWR VPWR _09314_/X sky130_fd_sc_hd__buf_1
XFILLER_34_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09245_ _09245_/A VGND VGND VPWR VPWR _09245_/X sky130_fd_sc_hd__buf_1
XFILLER_22_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09176_ _09176_/A VGND VGND VPWR VPWR _09176_/X sky130_fd_sc_hd__buf_1
XFILLER_135_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08127_ _08129_/A VGND VGND VPWR VPWR _08127_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08058_ _14312_/Q VGND VGND VPWR VPWR _08059_/A sky130_fd_sc_hd__buf_1
XFILLER_135_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10020_ _10389_/A VGND VGND VPWR VPWR _10020_/X sky130_fd_sc_hd__buf_1
XFILLER_49_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11971_ _11971_/A VGND VGND VPWR VPWR _11971_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13710_ _14973_/Q _15069_/Q _15037_/Q _15101_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13710_/X sky130_fd_sc_hd__mux4_2
X_10922_ _10922_/A VGND VGND VPWR VPWR _10929_/A sky130_fd_sc_hd__buf_1
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14690_ _10948_/X _14690_/D VGND VGND VPWR VPWR _14690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13641_ _13640_/X _07376_/Y _13641_/S VGND VGND VPWR VPWR _13641_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10853_ _10874_/A VGND VGND VPWR VPWR _10853_/X sky130_fd_sc_hd__buf_1
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _14096_/X _14101_/X _13648_/S VGND VGND VPWR VPWR _13572_/X sky130_fd_sc_hd__mux2_1
X_10784_ _10815_/A VGND VGND VPWR VPWR _10784_/X sky130_fd_sc_hd__buf_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15311_ _08469_/X _15311_/D VGND VGND VPWR VPWR _15311_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _15592_/Q VGND VGND VPWR VPWR _12524_/A sky130_fd_sc_hd__inv_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15242_ _08752_/X _15242_/D VGND VGND VPWR VPWR _15242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12454_ _12444_/Y _12449_/X _12453_/X VGND VGND VPWR VPWR _12454_/Y sky130_fd_sc_hd__o21ai_1
X_11405_ _11415_/A VGND VGND VPWR VPWR _11405_/X sky130_fd_sc_hd__buf_1
X_15173_ _09030_/X _15173_/D VGND VGND VPWR VPWR _15173_/Q sky130_fd_sc_hd__dfxtp_1
X_12385_ _13185_/X _12383_/X _12384_/X _12379_/Y VGND VGND VPWR VPWR _12385_/X sky130_fd_sc_hd__o22a_1
XFILLER_153_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14124_ _15187_/Q _15155_/Q _14771_/Q _14803_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14124_/X sky130_fd_sc_hd__mux4_1
X_11336_ _14591_/Q _11332_/X _11081_/X _11335_/X VGND VGND VPWR VPWR _14591_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14055_ _15130_/Q _15354_/Q _15322_/Q _15290_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14055_/X sky130_fd_sc_hd__mux4_1
X_11267_ _11269_/A VGND VGND VPWR VPWR _11267_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13006_ _14350_/Q VGND VGND VPWR VPWR _13006_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10218_ _10218_/A VGND VGND VPWR VPWR _10218_/X sky130_fd_sc_hd__buf_1
X_11198_ _11567_/A VGND VGND VPWR VPWR _11198_/X sky130_fd_sc_hd__buf_1
XFILLER_95_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10149_ _10167_/A VGND VGND VPWR VPWR _10149_/X sky130_fd_sc_hd__buf_1
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14957_ _09885_/X _14957_/D VGND VGND VPWR VPWR _14957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13908_ _14505_/Q _14473_/Q _14441_/Q _14409_/Q _13918_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13908_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14888_ _10162_/X _14888_/D VGND VGND VPWR VPWR _14888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13839_ _14832_/Q _14864_/Q _14896_/Q _14928_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13839_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07360_ _07362_/B VGND VGND VPWR VPWR _07360_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15509_ _15509_/CLK _15509_/D VGND VGND VPWR VPWR _15509_/Q sky130_fd_sc_hd__dfxtp_1
X_07291_ _07291_/A _13427_/X VGND VGND VPWR VPWR _15605_/D sky130_fd_sc_hd__and2_1
XFILLER_30_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09030_ _09030_/A VGND VGND VPWR VPWR _09030_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09932_ _14946_/Q _09927_/X _09928_/X _09931_/X VGND VGND VPWR VPWR _14946_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09863_ _09867_/A VGND VGND VPWR VPWR _09863_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08814_ _08827_/A VGND VGND VPWR VPWR _08814_/X sky130_fd_sc_hd__buf_1
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09794_ _09830_/A VGND VGND VPWR VPWR _09817_/A sky130_fd_sc_hd__buf_2
XFILLER_86_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08745_ _15245_/Q _08742_/X _08485_/X _08744_/X VGND VGND VPWR VPWR _15245_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_208 _13504_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08676_ _08676_/A VGND VGND VPWR VPWR _08676_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_219 _09205_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07627_ _07631_/A VGND VGND VPWR VPWR _07630_/A sky130_fd_sc_hd__buf_1
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07558_ _12986_/A VGND VGND VPWR VPWR _07558_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07489_ _07517_/A _13520_/X VGND VGND VPWR VPWR _15530_/D sky130_fd_sc_hd__and2_1
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09228_ _09228_/A VGND VGND VPWR VPWR _09228_/X sky130_fd_sc_hd__buf_1
XFILLER_10_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09159_ _09159_/A VGND VGND VPWR VPWR _09159_/X sky130_fd_sc_hd__buf_1
XFILLER_147_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12170_ _15542_/Q VGND VGND VPWR VPWR _12271_/A sky130_fd_sc_hd__inv_2
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11121_ _11489_/A VGND VGND VPWR VPWR _11121_/X sky130_fd_sc_hd__buf_1
XFILLER_150_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11052_ _11054_/A VGND VGND VPWR VPWR _11052_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10003_ _10371_/A VGND VGND VPWR VPWR _10003_/X sky130_fd_sc_hd__buf_1
XFILLER_49_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14811_ _10468_/X _14811_/D VGND VGND VPWR VPWR _14811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11954_ _11962_/A VGND VGND VPWR VPWR _11954_/X sky130_fd_sc_hd__clkbuf_1
X_14742_ _10730_/X _14742_/D VGND VGND VPWR VPWR _14742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10905_ _10905_/A VGND VGND VPWR VPWR _10905_/X sky130_fd_sc_hd__buf_1
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14673_ _11012_/X _14673_/D VGND VGND VPWR VPWR _14673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11885_ _11889_/A VGND VGND VPWR VPWR _11885_/X sky130_fd_sc_hd__clkbuf_1
X_13624_ _14226_/X _14231_/X _13648_/S VGND VGND VPWR VPWR _13624_/X sky130_fd_sc_hd__mux2_2
Xrepeater11 _15561_/Q VGND VGND VPWR VPWR _13418_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10836_ _10862_/A VGND VGND VPWR VPWR _10847_/A sky130_fd_sc_hd__buf_1
XFILLER_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater22 _13918_/S0 VGND VGND VPWR VPWR _13860_/S0 sky130_fd_sc_hd__clkbuf_16
Xrepeater33 _14398_/Q VGND VGND VPWR VPWR _14266_/S1 sky130_fd_sc_hd__clkbuf_16
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater44 _14238_/S0 VGND VGND VPWR VPWR _14180_/S0 sky130_fd_sc_hd__clkbuf_16
X_13555_ _13554_/X _13083_/X _14337_/Q VGND VGND VPWR VPWR _13555_/X sky130_fd_sc_hd__mux2_1
X_10767_ _10767_/A VGND VGND VPWR VPWR _10767_/X sky130_fd_sc_hd__buf_1
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12506_ _12498_/X _12347_/X _12495_/A _12505_/X VGND VGND VPWR VPWR _12507_/A sky130_fd_sc_hd__o22a_1
XFILLER_145_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13486_ _13485_/X rdata[12] _13516_/S VGND VGND VPWR VPWR _13486_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10698_ _11459_/A VGND VGND VPWR VPWR _10698_/X sky130_fd_sc_hd__buf_1
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15225_ _08824_/X _15225_/D VGND VGND VPWR VPWR _15225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12437_ _12437_/A VGND VGND VPWR VPWR _12505_/A sky130_fd_sc_hd__buf_1
XFILLER_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15156_ _09092_/X _15156_/D VGND VGND VPWR VPWR _15156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12368_ _12620_/A VGND VGND VPWR VPWR _12368_/X sky130_fd_sc_hd__buf_1
X_14107_ _14645_/Q _14613_/Q _14581_/Q _15381_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14107_/X sky130_fd_sc_hd__mux4_2
X_11319_ _11319_/A VGND VGND VPWR VPWR _11319_/X sky130_fd_sc_hd__buf_1
X_15087_ _09368_/X _15087_/D VGND VGND VPWR VPWR _15087_/Q sky130_fd_sc_hd__dfxtp_1
X_12299_ _15585_/Q VGND VGND VPWR VPWR _12330_/A sky130_fd_sc_hd__inv_2
XFILLER_113_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14038_ _14524_/Q _14492_/Q _14460_/Q _14428_/Q _14395_/Q _14060_/S1 VGND VGND VPWR
+ VPWR _14038_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08530_ _15302_/Q _08520_/X _08529_/X _08524_/X VGND VGND VPWR VPWR _15302_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08461_ _15313_/Q _08445_/X _08460_/X _08449_/X VGND VGND VPWR VPWR _15313_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07412_ _07416_/A VGND VGND VPWR VPWR _07415_/A sky130_fd_sc_hd__clkbuf_1
X_08392_ _15324_/Q _08387_/X _08390_/X _08391_/X VGND VGND VPWR VPWR _15324_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07343_ _07345_/B VGND VGND VPWR VPWR _07343_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07274_ _07274_/A VGND VGND VPWR VPWR _07283_/A sky130_fd_sc_hd__buf_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09013_ _15179_/Q _09006_/X _08887_/X _09008_/X VGND VGND VPWR VPWR _15179_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09915_ _09915_/A VGND VGND VPWR VPWR _09915_/X sky130_fd_sc_hd__buf_1
X_09846_ _09846_/A VGND VGND VPWR VPWR _09846_/X sky130_fd_sc_hd__buf_1
XFILLER_58_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09777_ _09797_/A VGND VGND VPWR VPWR _09777_/X sky130_fd_sc_hd__buf_1
XFILLER_27_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08728_ _15250_/Q _08723_/X _08454_/X _08724_/X VGND VGND VPWR VPWR _15250_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08659_ _08659_/A VGND VGND VPWR VPWR _08659_/X sky130_fd_sc_hd__clkbuf_1
X_11670_ _14504_/Q _11664_/X _11549_/X _11665_/X VGND VGND VPWR VPWR _14504_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10621_ _10625_/A VGND VGND VPWR VPWR _10621_/X sky130_fd_sc_hd__clkbuf_1
X_13340_ _13418_/X _13417_/X _13415_/S VGND VGND VPWR VPWR _13340_/X sky130_fd_sc_hd__mux2_1
X_10552_ _10565_/A VGND VGND VPWR VPWR _10553_/A sky130_fd_sc_hd__buf_1
XFILLER_6_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13271_ _12762_/X _12785_/A _13418_/S VGND VGND VPWR VPWR _13271_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10483_ _10514_/A VGND VGND VPWR VPWR _10505_/A sky130_fd_sc_hd__buf_2
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15010_ _09699_/X _15010_/D VGND VGND VPWR VPWR _15010_/Q sky130_fd_sc_hd__dfxtp_1
X_12222_ _15530_/Q VGND VGND VPWR VPWR _12223_/A sky130_fd_sc_hd__inv_2
X_12153_ _15543_/Q VGND VGND VPWR VPWR _12160_/A sky130_fd_sc_hd__inv_2
XFILLER_78_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11104_ _11471_/A VGND VGND VPWR VPWR _11104_/X sky130_fd_sc_hd__buf_1
XFILLER_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12084_ _12094_/A VGND VGND VPWR VPWR _12084_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11035_ _14667_/Q _11025_/X _10794_/X _11027_/X VGND VGND VPWR VPWR _14667_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12986_ _12986_/A _12993_/B VGND VGND VPWR VPWR _12986_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14725_ _10822_/X _14725_/D VGND VGND VPWR VPWR _14725_/Q sky130_fd_sc_hd__dfxtp_1
X_11937_ _11947_/A VGND VGND VPWR VPWR _11937_/X sky130_fd_sc_hd__buf_1
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11868_ _11868_/A VGND VGND VPWR VPWR _11868_/X sky130_fd_sc_hd__clkbuf_1
X_14656_ _11074_/X _14656_/D VGND VGND VPWR VPWR _14656_/Q sky130_fd_sc_hd__dfxtp_1
X_10819_ _11557_/A VGND VGND VPWR VPWR _10819_/X sky130_fd_sc_hd__buf_1
X_13607_ _13606_/X _13070_/X _14337_/Q VGND VGND VPWR VPWR _13607_/X sky130_fd_sc_hd__mux2_1
X_11799_ _11811_/A VGND VGND VPWR VPWR _11800_/A sky130_fd_sc_hd__buf_1
X_14587_ _11349_/X _14587_/D VGND VGND VPWR VPWR _14587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13538_ _13537_/X _14332_/D _15506_/Q VGND VGND VPWR VPWR _13538_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13469_ _13468_/X _13077_/X _14336_/Q VGND VGND VPWR VPWR _13469_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15208_ _08900_/X _15208_/D VGND VGND VPWR VPWR _15208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15139_ _09147_/X _15139_/D VGND VGND VPWR VPWR _15139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07961_ _07971_/A VGND VGND VPWR VPWR _07961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09700_ _09700_/A _11317_/B VGND VGND VPWR VPWR _09713_/A sky130_fd_sc_hd__or2_2
XFILLER_101_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07892_ _07891_/A _07891_/B _07882_/X _07891_/Y VGND VGND VPWR VPWR _15434_/D sky130_fd_sc_hd__o211a_1
XFILLER_95_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09631_ _10770_/A VGND VGND VPWR VPWR _10383_/A sky130_fd_sc_hd__buf_1
XFILLER_110_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09562_ _09577_/A VGND VGND VPWR VPWR _09562_/X sky130_fd_sc_hd__buf_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08513_ _08531_/A VGND VGND VPWR VPWR _08526_/A sky130_fd_sc_hd__buf_1
XFILLER_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09493_ _09495_/A VGND VGND VPWR VPWR _09493_/X sky130_fd_sc_hd__clkbuf_1
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08444_ _08451_/A VGND VGND VPWR VPWR _08444_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ _14331_/Q VGND VGND VPWR VPWR _10690_/A sky130_fd_sc_hd__buf_1
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07326_ _07329_/B VGND VGND VPWR VPWR _07326_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07257_ _07257_/A VGND VGND VPWR VPWR _07260_/A sky130_fd_sc_hd__buf_1
XFILLER_152_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07188_ _07235_/A VGND VGND VPWR VPWR _07188_/X sky130_fd_sc_hd__buf_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09829_ _14975_/Q _09825_/X _09546_/X _09828_/X VGND VGND VPWR VPWR _14975_/D sky130_fd_sc_hd__a22o_1
XFILLER_74_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12840_ _12838_/A _12261_/A _12839_/Y VGND VGND VPWR VPWR _12840_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12771_ _12875_/A VGND VGND VPWR VPWR _12929_/A sky130_fd_sc_hd__buf_1
XFILLER_27_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14510_ _11647_/X _14510_/D VGND VGND VPWR VPWR _14510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11722_ _11722_/A VGND VGND VPWR VPWR _11722_/X sky130_fd_sc_hd__buf_1
X_15490_ _15597_/CLK _15490_/D VGND VGND VPWR VPWR wdata[16] sky130_fd_sc_hd__dfxtp_2
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _11889_/X _14441_/D VGND VGND VPWR VPWR _14441_/Q sky130_fd_sc_hd__dfxtp_1
X_11653_ _11653_/A VGND VGND VPWR VPWR _11674_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _10606_/A VGND VGND VPWR VPWR _10604_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14372_ _14372_/CLK instruction[1] VGND VGND VPWR VPWR _14372_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11584_ _14529_/Q _11578_/X _11437_/X _11581_/X VGND VGND VPWR VPWR _14529_/D sky130_fd_sc_hd__a22o_1
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13323_ _12211_/X _12875_/B _15561_/Q VGND VGND VPWR VPWR _13323_/X sky130_fd_sc_hd__mux2_1
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10535_ _10535_/A VGND VGND VPWR VPWR _10535_/X sky130_fd_sc_hd__buf_1
XFILLER_10_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13254_ _13312_/X _13311_/X _13393_/S VGND VGND VPWR VPWR _13254_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10466_ _10475_/A VGND VGND VPWR VPWR _10466_/X sky130_fd_sc_hd__buf_1
XFILLER_142_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12205_ _15570_/Q VGND VGND VPWR VPWR _12779_/A sky130_fd_sc_hd__inv_2
X_13185_ _13184_/X _13268_/X _15565_/Q VGND VGND VPWR VPWR _13185_/X sky130_fd_sc_hd__mux2_1
X_10397_ _14829_/Q _10393_/X _10394_/X _10396_/X VGND VGND VPWR VPWR _14829_/D sky130_fd_sc_hd__a22o_1
X_12136_ _15546_/Q VGND VGND VPWR VPWR _12142_/A sky130_fd_sc_hd__inv_2
XFILLER_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12067_ _12071_/A VGND VGND VPWR VPWR _12156_/A sky130_fd_sc_hd__buf_1
X_11018_ _11018_/A VGND VGND VPWR VPWR _11023_/A sky130_fd_sc_hd__buf_1
XFILLER_38_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12969_ _12600_/X _12955_/Y _12706_/A _12967_/X _12968_/X VGND VGND VPWR VPWR _12969_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14708_ _10890_/X _14708_/D VGND VGND VPWR VPWR _14708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14639_ _11151_/X _14639_/D VGND VGND VPWR VPWR _14639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08160_ _15380_/Q _08153_/X _08011_/X _08155_/X VGND VGND VPWR VPWR _15380_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07111_ rst VGND VGND VPWR VPWR _07182_/A sky130_fd_sc_hd__inv_2
X_08091_ _08091_/A VGND VGND VPWR VPWR _08091_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08993_ _08993_/A VGND VGND VPWR VPWR _08993_/X sky130_fd_sc_hd__buf_1
XFILLER_114_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07944_ _07944_/A VGND VGND VPWR VPWR _07944_/X sky130_fd_sc_hd__buf_1
XFILLER_96_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07875_ _07875_/A VGND VGND VPWR VPWR _07884_/B sky130_fd_sc_hd__buf_1
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09614_ _15027_/Q _09610_/X _09612_/X _09613_/X VGND VGND VPWR VPWR _15027_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09545_ _10683_/A VGND VGND VPWR VPWR _10314_/A sky130_fd_sc_hd__buf_1
XFILLER_37_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09476_ _09476_/A VGND VGND VPWR VPWR _09476_/X sky130_fd_sc_hd__buf_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08427_ _09211_/A VGND VGND VPWR VPWR _08427_/X sky130_fd_sc_hd__buf_1
XFILLER_12_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ _08374_/A VGND VGND VPWR VPWR _08358_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07309_ _07298_/X _07301_/X _07559_/D _07321_/C _07308_/X VGND VGND VPWR VPWR _07314_/A
+ sky130_fd_sc_hd__o221a_2
X_08289_ _15345_/Q _08282_/X _08026_/X _08283_/X VGND VGND VPWR VPWR _15345_/D sky130_fd_sc_hd__a22o_1
X_10320_ _10320_/A VGND VGND VPWR VPWR _10320_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10251_ _10255_/A VGND VGND VPWR VPWR _10251_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10182_ _10194_/A VGND VGND VPWR VPWR _10183_/A sky130_fd_sc_hd__buf_1
XFILLER_105_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14990_ _09772_/X _14990_/D VGND VGND VPWR VPWR _14990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13941_ _13937_/X _13938_/X _13939_/X _13940_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13941_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13872_ _15212_/Q _14540_/Q _14988_/Q _15404_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13872_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15611_ _15648_/CLK _15611_/D VGND VGND VPWR VPWR pc[6] sky130_fd_sc_hd__dfxtp_1
X_12823_ _12823_/A _12883_/A VGND VGND VPWR VPWR _12824_/A sky130_fd_sc_hd__or2_1
XFILLER_15_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15542_ _15621_/CLK _15542_/D VGND VGND VPWR VPWR _15542_/Q sky130_fd_sc_hd__dfxtp_1
X_12754_ _12754_/A VGND VGND VPWR VPWR _12758_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11705_ _11723_/A VGND VGND VPWR VPWR _11705_/X sky130_fd_sc_hd__buf_1
X_15473_ _15599_/CLK _15473_/D VGND VGND VPWR VPWR _15473_/Q sky130_fd_sc_hd__dfxtp_1
X_12685_ _12685_/A VGND VGND VPWR VPWR _12735_/A sky130_fd_sc_hd__clkbuf_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ _11638_/A VGND VGND VPWR VPWR _11636_/X sky130_fd_sc_hd__clkbuf_1
X_14424_ _11949_/X _14424_/D VGND VGND VPWR VPWR _14424_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14355_ _15652_/CLK pc[16] VGND VGND VPWR VPWR _14355_/Q sky130_fd_sc_hd__dfxtp_1
X_11567_ _11567_/A VGND VGND VPWR VPWR _11567_/X sky130_fd_sc_hd__buf_1
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13306_ _12847_/A _12838_/X _15561_/Q VGND VGND VPWR VPWR _13306_/X sky130_fd_sc_hd__mux2_1
X_10518_ _14797_/Q _10515_/X _10394_/X _10517_/X VGND VGND VPWR VPWR _14797_/D sky130_fd_sc_hd__a22o_1
X_14286_ _14282_/X _14283_/X _14284_/X _14285_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14286_/X sky130_fd_sc_hd__mux4_2
XFILLER_143_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11498_ _11498_/A VGND VGND VPWR VPWR _11498_/X sky130_fd_sc_hd__buf_1
X_13237_ _12662_/X _12703_/A _13418_/S VGND VGND VPWR VPWR _13237_/X sky130_fd_sc_hd__mux2_1
X_10449_ _10449_/A VGND VGND VPWR VPWR _10460_/A sky130_fd_sc_hd__buf_1
XFILLER_124_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13168_ _13172_/X _13182_/X _15562_/Q VGND VGND VPWR VPWR _13168_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12119_ _15547_/Q VGND VGND VPWR VPWR _12635_/A sky130_fd_sc_hd__inv_2
X_13099_ _15645_/Q data_address[10] _15667_/Q VGND VGND VPWR VPWR _13099_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07660_ _07660_/A VGND VGND VPWR VPWR _07660_/X sky130_fd_sc_hd__buf_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07591_ _07591_/A _13074_/X VGND VGND VPWR VPWR _15489_/D sky130_fd_sc_hd__and2_1
XFILLER_19_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09330_ _15099_/Q _09326_/X _09188_/X _09327_/X VGND VGND VPWR VPWR _15099_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09261_ _09266_/A VGND VGND VPWR VPWR _09261_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08212_ _08216_/A VGND VGND VPWR VPWR _08212_/X sky130_fd_sc_hd__clkbuf_1
X_09192_ _09192_/A VGND VGND VPWR VPWR _09192_/X sky130_fd_sc_hd__buf_1
XFILLER_119_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08143_ _08143_/A VGND VGND VPWR VPWR _08143_/X sky130_fd_sc_hd__buf_1
X_08074_ _08074_/A VGND VGND VPWR VPWR _08074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08976_ _08994_/A VGND VGND VPWR VPWR _08976_/X sky130_fd_sc_hd__buf_1
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07927_ _07927_/A VGND VGND VPWR VPWR _07927_/X sky130_fd_sc_hd__buf_1
X_07858_ _07863_/A _07863_/B VGND VGND VPWR VPWR _07864_/B sky130_fd_sc_hd__or2_1
XFILLER_45_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07789_ _07789_/A _07789_/B VGND VGND VPWR VPWR _07789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09528_ _09542_/A VGND VGND VPWR VPWR _09547_/A sky130_fd_sc_hd__inv_2
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09459_ _15062_/Q _09456_/X _09211_/X _09458_/X VGND VGND VPWR VPWR _15062_/D sky130_fd_sc_hd__a22o_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12470_ _15558_/Q VGND VGND VPWR VPWR _12470_/X sky130_fd_sc_hd__buf_1
XFILLER_12_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11421_ _14565_/Q _11414_/X _11195_/X _11415_/X VGND VGND VPWR VPWR _14565_/D sky130_fd_sc_hd__a22o_1
XFILLER_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14140_ _14962_/Q _15058_/Q _15026_/Q _15090_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14140_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11352_ _14586_/Q _11343_/X _11104_/X _11344_/X VGND VGND VPWR VPWR _14586_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10303_ _10303_/A VGND VGND VPWR VPWR _10303_/X sky130_fd_sc_hd__buf_1
XFILLER_152_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14071_ _14067_/X _14068_/X _14069_/X _14070_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14071_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11283_ _11283_/A VGND VGND VPWR VPWR _11303_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13022_ _14366_/Q VGND VGND VPWR VPWR _13022_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10234_ _10236_/A VGND VGND VPWR VPWR _10234_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10165_ _10171_/A VGND VGND VPWR VPWR _10165_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14973_ _09834_/X _14973_/D VGND VGND VPWR VPWR _14973_/Q sky130_fd_sc_hd__dfxtp_1
X_10096_ _10102_/A VGND VGND VPWR VPWR _10096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13924_ _15175_/Q _15143_/Q _14759_/Q _14791_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13924_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13855_ _15118_/Q _15342_/Q _15310_/Q _15278_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13855_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12806_ _12806_/A VGND VGND VPWR VPWR _12812_/A sky130_fd_sc_hd__buf_4
XFILLER_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13786_ _13782_/X _13783_/X _13784_/X _13785_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13786_/X sky130_fd_sc_hd__mux4_2
X_10998_ _14678_/Q _10995_/X _10734_/X _10997_/X VGND VGND VPWR VPWR _14678_/D sky130_fd_sc_hd__a22o_1
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15525_ _15597_/CLK _15525_/D VGND VGND VPWR VPWR _15525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12737_ _12737_/A _12737_/B VGND VGND VPWR VPWR _12913_/B sky130_fd_sc_hd__nor2_2
XFILLER_31_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15456_ _15456_/CLK _15456_/D VGND VGND VPWR VPWR data_address[29] sky130_fd_sc_hd__dfxtp_4
X_12668_ _12668_/A VGND VGND VPWR VPWR _12668_/X sky130_fd_sc_hd__buf_1
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _12004_/X _14407_/D VGND VGND VPWR VPWR _14407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11619_ _11619_/A VGND VGND VPWR VPWR _11628_/A sky130_fd_sc_hd__buf_1
X_15387_ _08137_/X _15387_/D VGND VGND VPWR VPWR _15387_/Q sky130_fd_sc_hd__dfxtp_1
X_12599_ _12599_/A VGND VGND VPWR VPWR _12599_/X sky130_fd_sc_hd__buf_1
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14338_ _12017_/X _15670_/Q VGND VGND VPWR VPWR _14338_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14269_ _14821_/Q _14853_/Q _14885_/Q _14917_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14269_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08830_ _09200_/A VGND VGND VPWR VPWR _08830_/X sky130_fd_sc_hd__buf_1
XFILLER_39_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08761_ _08761_/A VGND VGND VPWR VPWR _08761_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07712_ _07706_/A _07711_/X _07687_/A _13137_/X VGND VGND VPWR VPWR _07712_/X sky130_fd_sc_hd__o22a_1
XFILLER_38_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08692_ _08692_/A VGND VGND VPWR VPWR _08692_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07643_ _15604_/Q VGND VGND VPWR VPWR _07660_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07574_ _07582_/A VGND VGND VPWR VPWR _07577_/A sky130_fd_sc_hd__buf_1
XFILLER_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09313_ _09376_/A VGND VGND VPWR VPWR _09336_/A sky130_fd_sc_hd__buf_2
XFILLER_22_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09244_ _09254_/A VGND VGND VPWR VPWR _09244_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09175_ _09175_/A VGND VGND VPWR VPWR _09175_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08126_ _15391_/Q _08122_/X _07951_/X _08125_/X VGND VGND VPWR VPWR _15391_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08057_ _08067_/A VGND VGND VPWR VPWR _08057_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08959_ _08959_/A VGND VGND VPWR VPWR _08959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11970_ _14418_/Q _11966_/X _08021_/A _11967_/X VGND VGND VPWR VPWR _14418_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10921_ _14699_/Q _10914_/X _10794_/X _10916_/X VGND VGND VPWR VPWR _14699_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10852_ _10913_/A VGND VGND VPWR VPWR _10874_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13640_ _14266_/X _14271_/X _13648_/S VGND VGND VPWR VPWR _13640_/X sky130_fd_sc_hd__mux2_2
XFILLER_112_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10783_ _10783_/A VGND VGND VPWR VPWR _10815_/A sky130_fd_sc_hd__buf_1
X_13571_ _13570_/X _13079_/X _14337_/Q VGND VGND VPWR VPWR _13571_/X sky130_fd_sc_hd__mux2_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_clk _14315_/CLK VGND VGND VPWR VPWR _15662_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15310_ _08475_/X _15310_/D VGND VGND VPWR VPWR _15310_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _12522_/A VGND VGND VPWR VPWR _12522_/X sky130_fd_sc_hd__buf_1
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15241_ _08757_/X _15241_/D VGND VGND VPWR VPWR _15241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12453_ _12450_/X _12447_/A _13176_/X _12451_/X _12452_/X VGND VGND VPWR VPWR _12453_/X
+ sky130_fd_sc_hd__o221a_1
X_11404_ _11414_/A VGND VGND VPWR VPWR _11404_/X sky130_fd_sc_hd__buf_1
X_12384_ _12448_/A VGND VGND VPWR VPWR _12384_/X sky130_fd_sc_hd__buf_1
X_15172_ _09034_/X _15172_/D VGND VGND VPWR VPWR _15172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14123_ _14675_/Q _15251_/Q _14739_/Q _14707_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14123_/X sky130_fd_sc_hd__mux4_2
X_11335_ _11355_/A VGND VGND VPWR VPWR _11335_/X sky130_fd_sc_hd__buf_1
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11266_ _14611_/Q _11264_/X _11134_/X _11265_/X VGND VGND VPWR VPWR _14611_/D sky130_fd_sc_hd__a22o_1
X_14054_ _15194_/Q _15162_/Q _14778_/Q _14810_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14054_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13005_ _14349_/Q VGND VGND VPWR VPWR _13005_/Y sky130_fd_sc_hd__inv_2
X_10217_ _10217_/A VGND VGND VPWR VPWR _10217_/X sky130_fd_sc_hd__buf_1
X_11197_ _11200_/A VGND VGND VPWR VPWR _11197_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10148_ _10148_/A VGND VGND VPWR VPWR _10167_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10079_ _14912_/Q _10071_/X _09938_/X _10074_/X VGND VGND VPWR VPWR _14912_/D sky130_fd_sc_hd__a22o_1
X_14956_ _09893_/X _14956_/D VGND VGND VPWR VPWR _14956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13907_ _14633_/Q _14601_/Q _14569_/Q _15369_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13907_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14887_ _10165_/X _14887_/D VGND VGND VPWR VPWR _14887_/Q sky130_fd_sc_hd__dfxtp_1
X_13838_ _14512_/Q _14480_/Q _14448_/Q _14416_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13838_/X sky130_fd_sc_hd__mux4_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13769_ _14839_/Q _14871_/Q _14903_/Q _14935_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13769_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_42_clk clkbuf_opt_7_clk/X VGND VGND VPWR VPWR _15527_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15508_ _15599_/CLK _15508_/D VGND VGND VPWR VPWR _15508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07290_ _07291_/A _13426_/X VGND VGND VPWR VPWR _15606_/D sky130_fd_sc_hd__and2_1
XFILLER_30_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15439_ _15621_/CLK _15439_/D VGND VGND VPWR VPWR data_address[12] sky130_fd_sc_hd__dfxtp_4
XFILLER_116_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09931_ _09931_/A VGND VGND VPWR VPWR _09931_/X sky130_fd_sc_hd__buf_1
X_09862_ _09880_/A VGND VGND VPWR VPWR _09867_/A sky130_fd_sc_hd__buf_1
XFILLER_86_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08813_ _09184_/A VGND VGND VPWR VPWR _08813_/X sky130_fd_sc_hd__buf_1
XFILLER_85_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09793_ _14984_/Q _09787_/X _09672_/X _09788_/X VGND VGND VPWR VPWR _14984_/D sky130_fd_sc_hd__a22o_1
X_08744_ _08763_/A VGND VGND VPWR VPWR _08744_/X sky130_fd_sc_hd__buf_1
XFILLER_66_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_209 _13501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08675_ _15264_/Q _08666_/X _08361_/X _08669_/X VGND VGND VPWR VPWR _15264_/D sky130_fd_sc_hd__a22o_1
X_07626_ _07626_/A _12984_/C VGND VGND VPWR VPWR _15471_/D sky130_fd_sc_hd__nor2_1
X_07557_ _12986_/A _12993_/A _07297_/A VGND VGND VPWR VPWR _07557_/X sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_33_clk _14315_/CLK VGND VGND VPWR VPWR _15667_/CLK sky130_fd_sc_hd__clkbuf_16
X_07488_ _07569_/A VGND VGND VPWR VPWR _07517_/A sky130_fd_sc_hd__buf_1
XFILLER_22_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09227_ _09227_/A VGND VGND VPWR VPWR _09227_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09158_ _09158_/A VGND VGND VPWR VPWR _09158_/X sky130_fd_sc_hd__clkbuf_1
X_08109_ _08109_/A VGND VGND VPWR VPWR _08109_/X sky130_fd_sc_hd__buf_1
X_09089_ _09089_/A VGND VGND VPWR VPWR _09094_/A sky130_fd_sc_hd__buf_1
XFILLER_107_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11120_ _11147_/A VGND VGND VPWR VPWR _11120_/X sky130_fd_sc_hd__buf_1
XFILLER_122_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11051_ _14662_/Q _11046_/X _10819_/X _11047_/X VGND VGND VPWR VPWR _14662_/D sky130_fd_sc_hd__a22o_1
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10002_ _10002_/A VGND VGND VPWR VPWR _10002_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14810_ _10470_/X _14810_/D VGND VGND VPWR VPWR _14810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14741_ _10738_/X _14741_/D VGND VGND VPWR VPWR _14741_/Q sky130_fd_sc_hd__dfxtp_1
X_11953_ _11964_/A VGND VGND VPWR VPWR _11962_/A sky130_fd_sc_hd__buf_1
XFILLER_44_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10904_ _10904_/A VGND VGND VPWR VPWR _10904_/X sky130_fd_sc_hd__buf_1
XFILLER_60_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14672_ _11014_/X _14672_/D VGND VGND VPWR VPWR _14672_/Q sky130_fd_sc_hd__dfxtp_1
X_11884_ _14443_/Q _11875_/X _08059_/A _11877_/X VGND VGND VPWR VPWR _14443_/D sky130_fd_sc_hd__a22o_1
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13623_ _13622_/X _13066_/X _14337_/Q VGND VGND VPWR VPWR _13623_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR _14328_/CLK sky130_fd_sc_hd__clkbuf_1
X_10835_ _10901_/A VGND VGND VPWR VPWR _10862_/A sky130_fd_sc_hd__buf_2
XFILLER_13_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater12 _13946_/S1 VGND VGND VPWR VPWR _13966_/S1 sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_24_clk _14397_/CLK VGND VGND VPWR VPWR _14385_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater23 _13918_/S0 VGND VGND VPWR VPWR _13825_/S0 sky130_fd_sc_hd__clkbuf_16
Xrepeater34 _14266_/S0 VGND VGND VPWR VPWR _14286_/S0 sky130_fd_sc_hd__clkbuf_16
Xrepeater45 _14238_/S0 VGND VGND VPWR VPWR _14145_/S0 sky130_fd_sc_hd__clkbuf_16
X_13554_ _13553_/X _14328_/D _15506_/Q VGND VGND VPWR VPWR _13554_/X sky130_fd_sc_hd__mux2_2
XFILLER_9_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10766_ _11514_/A VGND VGND VPWR VPWR _10766_/X sky130_fd_sc_hd__buf_1
XFILLER_13_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12505_ _12505_/A VGND VGND VPWR VPWR _12505_/X sky130_fd_sc_hd__buf_1
X_13485_ _13846_/X _13851_/X _13521_/S VGND VGND VPWR VPWR _13485_/X sky130_fd_sc_hd__mux2_2
X_10697_ _10697_/A VGND VGND VPWR VPWR _11459_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15224_ _08829_/X _15224_/D VGND VGND VPWR VPWR _15224_/Q sky130_fd_sc_hd__dfxtp_1
X_12436_ _15589_/Q VGND VGND VPWR VPWR _12902_/A sky130_fd_sc_hd__inv_2
XFILLER_66_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15155_ _09094_/X _15155_/D VGND VGND VPWR VPWR _15155_/Q sky130_fd_sc_hd__dfxtp_1
X_12367_ _12367_/A VGND VGND VPWR VPWR _12620_/A sky130_fd_sc_hd__buf_1
XFILLER_153_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14106_ _14102_/X _14103_/X _14104_/X _14105_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14106_/X sky130_fd_sc_hd__mux4_2
X_11318_ _11330_/A VGND VGND VPWR VPWR _11319_/A sky130_fd_sc_hd__buf_1
X_15086_ _09370_/X _15086_/D VGND VGND VPWR VPWR _15086_/Q sky130_fd_sc_hd__dfxtp_1
X_12298_ _12346_/A VGND VGND VPWR VPWR _12298_/X sky130_fd_sc_hd__buf_1
XFILLER_141_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11249_ _11439_/A VGND VGND VPWR VPWR _11310_/A sky130_fd_sc_hd__buf_1
X_14037_ _14652_/Q _14620_/Q _14588_/Q _15388_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14037_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14939_ _09961_/X _14939_/D VGND VGND VPWR VPWR _14939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08460_ _09232_/A VGND VGND VPWR VPWR _08460_/X sky130_fd_sc_hd__buf_1
XFILLER_63_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07411_ _07411_/A _13567_/X VGND VGND VPWR VPWR _15582_/D sky130_fd_sc_hd__and2_1
XFILLER_35_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08391_ _08409_/A VGND VGND VPWR VPWR _08391_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_15_clk _14328_/CLK VGND VGND VPWR VPWR _15502_/CLK sky130_fd_sc_hd__clkbuf_16
X_07342_ _07494_/B _07339_/X _07495_/B _07341_/X VGND VGND VPWR VPWR _07345_/B sky130_fd_sc_hd__o22a_1
XFILLER_148_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07273_ _07273_/A _07273_/B VGND VGND VPWR VPWR _15619_/D sky130_fd_sc_hd__nor2_1
X_09012_ _09012_/A VGND VGND VPWR VPWR _09012_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09914_ _14949_/Q _09907_/X _09687_/X _09908_/X VGND VGND VPWR VPWR _14949_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09845_ _09845_/A VGND VGND VPWR VPWR _09845_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09776_ _09776_/A VGND VGND VPWR VPWR _09797_/A sky130_fd_sc_hd__buf_1
XFILLER_73_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08727_ _08731_/A VGND VGND VPWR VPWR _08727_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08658_ _15267_/Q _08552_/A _08545_/X _08555_/A VGND VGND VPWR VPWR _15267_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07609_ _07609_/A VGND VGND VPWR VPWR _07638_/A sky130_fd_sc_hd__buf_1
XFILLER_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08589_ _15289_/Q _08587_/X _08408_/X _08588_/X VGND VGND VPWR VPWR _15289_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10620_ _10640_/A VGND VGND VPWR VPWR _10625_/A sky130_fd_sc_hd__buf_2
XFILLER_139_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10551_ _10562_/A VGND VGND VPWR VPWR _10565_/A sky130_fd_sc_hd__inv_2
XFILLER_139_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13270_ _13271_/X _13283_/X _13415_/S VGND VGND VPWR VPWR _13270_/X sky130_fd_sc_hd__mux2_1
X_10482_ _10490_/A VGND VGND VPWR VPWR _10482_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12221_ _12862_/A _12220_/A _15531_/Q _12220_/Y VGND VGND VPWR VPWR _12863_/A sky130_fd_sc_hd__o22a_1
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12152_ _12692_/A _12151_/B _12151_/Y VGND VGND VPWR VPWR _12162_/A sky130_fd_sc_hd__a21oi_4
XFILLER_135_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11103_ _11111_/A VGND VGND VPWR VPWR _11103_/X sky130_fd_sc_hd__buf_1
X_12083_ _15584_/Q VGND VGND VPWR VPWR _12591_/A sky130_fd_sc_hd__inv_2
XFILLER_104_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11034_ _11036_/A VGND VGND VPWR VPWR _11034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12985_ _15506_/D VGND VGND VPWR VPWR _12993_/B sky130_fd_sc_hd__inv_2
XFILLER_80_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14724_ _10826_/X _14724_/D VGND VGND VPWR VPWR _14724_/Q sky130_fd_sc_hd__dfxtp_1
X_11936_ _11946_/A VGND VGND VPWR VPWR _11936_/X sky130_fd_sc_hd__buf_1
XFILLER_91_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14655_ _11077_/X _14655_/D VGND VGND VPWR VPWR _14655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11867_ _14448_/Q _11865_/X _08031_/A _11866_/X VGND VGND VPWR VPWR _14448_/D sky130_fd_sc_hd__a22o_1
X_13606_ _13605_/X _14315_/D _15506_/Q VGND VGND VPWR VPWR _13606_/X sky130_fd_sc_hd__mux2_1
X_10818_ _10818_/A VGND VGND VPWR VPWR _11557_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14586_ _11351_/X _14586_/D VGND VGND VPWR VPWR _14586_/Q sky130_fd_sc_hd__dfxtp_1
X_11798_ _11798_/A _11798_/B VGND VGND VPWR VPWR _11811_/A sky130_fd_sc_hd__or2_2
XFILLER_41_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13537_ _13536_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13537_/X sky130_fd_sc_hd__mux2_1
X_10749_ _10764_/A VGND VGND VPWR VPWR _10749_/X sky130_fd_sc_hd__buf_1
XFILLER_146_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13468_ _13467_/X rdata[18] _14338_/Q VGND VGND VPWR VPWR _13468_/X sky130_fd_sc_hd__mux2_1
X_15207_ _08903_/X _15207_/D VGND VGND VPWR VPWR _15207_/Q sky130_fd_sc_hd__dfxtp_1
X_12419_ _12403_/X _12412_/A _12414_/X _12415_/A VGND VGND VPWR VPWR _12904_/D sky130_fd_sc_hd__o22a_1
X_13399_ _12388_/X _12415_/X _13418_/S VGND VGND VPWR VPWR _13399_/X sky130_fd_sc_hd__mux2_1
X_15138_ _09149_/X _15138_/D VGND VGND VPWR VPWR _15138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15069_ _09433_/X _15069_/D VGND VGND VPWR VPWR _15069_/Q sky130_fd_sc_hd__dfxtp_1
X_07960_ _07975_/A VGND VGND VPWR VPWR _07971_/A sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_4_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR _14381_/CLK sky130_fd_sc_hd__clkbuf_16
X_07891_ _07891_/A _07891_/B VGND VGND VPWR VPWR _07891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09630_ _09630_/A VGND VGND VPWR VPWR _09630_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09561_ _09567_/A VGND VGND VPWR VPWR _09561_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08512_ _15305_/Q _08502_/X _08511_/X _08506_/X VGND VGND VPWR VPWR _15305_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09492_ _15052_/Q _09486_/X _09255_/X _09488_/X VGND VGND VPWR VPWR _15052_/D sky130_fd_sc_hd__a22o_1
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08443_ _15316_/Q _08424_/X _08442_/X _08429_/X VGND VGND VPWR VPWR _15316_/D sky130_fd_sc_hd__a22o_1
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ _08374_/A VGND VGND VPWR VPWR _08374_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07325_ _07512_/B _07319_/X _07491_/B _07324_/X VGND VGND VPWR VPWR _07329_/B sky130_fd_sc_hd__o22a_1
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07256_ _07256_/A _07256_/B VGND VGND VPWR VPWR _15631_/D sky130_fd_sc_hd__nor2_1
XFILLER_137_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07187_ _07247_/A VGND VGND VPWR VPWR _07235_/A sky130_fd_sc_hd__buf_1
XFILLER_117_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09828_ _09847_/A VGND VGND VPWR VPWR _09828_/X sky130_fd_sc_hd__buf_1
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09759_ _09761_/A VGND VGND VPWR VPWR _09759_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12770_ _12770_/A _13322_/X VGND VGND VPWR VPWR _12860_/B sky130_fd_sc_hd__or2_1
XFILLER_82_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11721_ _11721_/A VGND VGND VPWR VPWR _11721_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14440_ _11892_/X _14440_/D VGND VGND VPWR VPWR _14440_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11673_/A VGND VGND VPWR VPWR _11652_/X sky130_fd_sc_hd__buf_1
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ _14773_/Q _10597_/X _10359_/X _10599_/X VGND VGND VPWR VPWR _14773_/D sky130_fd_sc_hd__a22o_1
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ _14395_/CLK instruction[0] VGND VGND VPWR VPWR _14371_/Q sky130_fd_sc_hd__dfxtp_4
X_11583_ _11585_/A VGND VGND VPWR VPWR _11583_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13322_ _13323_/X _13355_/X _15562_/Q VGND VGND VPWR VPWR _13322_/X sky130_fd_sc_hd__mux2_1
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10534_ _10540_/A VGND VGND VPWR VPWR _10534_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13253_ _12730_/A _12737_/A _13418_/S VGND VGND VPWR VPWR _13253_/X sky130_fd_sc_hd__mux2_1
X_10465_ _10474_/A VGND VGND VPWR VPWR _10465_/X sky130_fd_sc_hd__buf_1
XFILLER_124_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12204_ _15570_/Q VGND VGND VPWR VPWR _12204_/X sky130_fd_sc_hd__buf_1
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13184_ _13183_/X _13225_/X _13393_/S VGND VGND VPWR VPWR _13184_/X sky130_fd_sc_hd__mux2_1
X_10396_ _10420_/A VGND VGND VPWR VPWR _10396_/X sky130_fd_sc_hd__buf_1
XFILLER_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12135_ _12135_/A VGND VGND VPWR VPWR _12144_/B sky130_fd_sc_hd__inv_2
XFILLER_97_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12066_ _12024_/A _12027_/A _13386_/X _12031_/A VGND VGND VPWR VPWR _12071_/A sky130_fd_sc_hd__o22a_1
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11017_ _14672_/Q _11015_/X _10766_/X _11016_/X VGND VGND VPWR VPWR _14672_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12968_ _13419_/X _12974_/B _07123_/A _13392_/X _12782_/A VGND VGND VPWR VPWR _12968_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_64_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14707_ _10893_/X _14707_/D VGND VGND VPWR VPWR _14707_/Q sky130_fd_sc_hd__dfxtp_1
X_11919_ _11919_/A VGND VGND VPWR VPWR _11919_/X sky130_fd_sc_hd__clkbuf_1
X_12899_ _12020_/X _12330_/X _12904_/C _12362_/X _12359_/X VGND VGND VPWR VPWR _12899_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_61_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14638_ _11155_/X _14638_/D VGND VGND VPWR VPWR _14638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14569_ _11409_/X _14569_/D VGND VGND VPWR VPWR _14569_/Q sky130_fd_sc_hd__dfxtp_1
X_07110_ _07893_/A VGND VGND VPWR VPWR _07909_/C sky130_fd_sc_hd__buf_1
XFILLER_118_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08090_ _14306_/Q VGND VGND VPWR VPWR _08091_/A sky130_fd_sc_hd__buf_1
XFILLER_118_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08992_ _08998_/A VGND VGND VPWR VPWR _08992_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07943_ _14333_/Q VGND VGND VPWR VPWR _07944_/A sky130_fd_sc_hd__buf_1
X_07874_ _07874_/A VGND VGND VPWR VPWR _07874_/X sky130_fd_sc_hd__buf_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09613_ _09628_/A VGND VGND VPWR VPWR _09613_/X sky130_fd_sc_hd__buf_1
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09544_ _09577_/A VGND VGND VPWR VPWR _09544_/X sky130_fd_sc_hd__buf_1
XFILLER_71_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09475_ _09475_/A VGND VGND VPWR VPWR _09475_/X sky130_fd_sc_hd__buf_1
XFILLER_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08426_ _10733_/A VGND VGND VPWR VPWR _09211_/A sky130_fd_sc_hd__buf_1
XFILLER_24_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08357_ _08357_/A VGND VGND VPWR VPWR _08374_/A sky130_fd_sc_hd__buf_2
XFILLER_137_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07308_ _07373_/A VGND VGND VPWR VPWR _07308_/X sky130_fd_sc_hd__buf_1
X_08288_ _08290_/A VGND VGND VPWR VPWR _08288_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07239_ _07288_/A _07239_/B _07239_/C VGND VGND VPWR VPWR _15640_/D sky130_fd_sc_hd__nor3_1
XFILLER_118_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10250_ _10261_/A VGND VGND VPWR VPWR _10255_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10181_ _11686_/A _10181_/B VGND VGND VPWR VPWR _10194_/A sky130_fd_sc_hd__or2_2
XFILLER_105_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13940_ _14950_/Q _15046_/Q _15014_/Q _15078_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13940_/X sky130_fd_sc_hd__mux4_2
XFILLER_115_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13871_ _13867_/X _13868_/X _13869_/X _13870_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13871_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15610_ _15666_/CLK _15610_/D VGND VGND VPWR VPWR pc[5] sky130_fd_sc_hd__dfxtp_1
X_12822_ _12878_/A VGND VGND VPWR VPWR _12883_/A sky130_fd_sc_hd__buf_1
XFILLER_28_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15541_ _15621_/CLK _15541_/D VGND VGND VPWR VPWR _15541_/Q sky130_fd_sc_hd__dfxtp_1
X_12753_ _12753_/A VGND VGND VPWR VPWR _12753_/X sky130_fd_sc_hd__buf_1
X_11704_ _11765_/A VGND VGND VPWR VPWR _11723_/A sky130_fd_sc_hd__buf_2
X_15472_ _15599_/CLK _15472_/D VGND VGND VPWR VPWR _15472_/Q sky130_fd_sc_hd__dfxtp_1
X_12684_ _12684_/A VGND VGND VPWR VPWR _12684_/X sky130_fd_sc_hd__buf_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _11951_/X _14423_/D VGND VGND VPWR VPWR _14423_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _14515_/Q _11633_/X _11502_/X _11634_/X VGND VGND VPWR VPWR _14515_/D sky130_fd_sc_hd__a22o_1
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14354_ _15621_/CLK pc[15] VGND VGND VPWR VPWR _14354_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _11569_/A VGND VGND VPWR VPWR _11566_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13305_ _13306_/X _13323_/X _15562_/Q VGND VGND VPWR VPWR _13305_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10517_ _10536_/A VGND VGND VPWR VPWR _10517_/X sky130_fd_sc_hd__buf_1
XFILLER_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14285_ _15107_/Q _15331_/Q _15299_/Q _15267_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14285_/X sky130_fd_sc_hd__mux4_1
X_11497_ _11505_/A VGND VGND VPWR VPWR _11497_/X sky130_fd_sc_hd__buf_1
XFILLER_115_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13236_ _13237_/X _13247_/X _13415_/S VGND VGND VPWR VPWR _13236_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10448_ _14816_/Q _10440_/X _10308_/X _10443_/X VGND VGND VPWR VPWR _14816_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13167_ _13166_/X _13244_/X _15565_/Q VGND VGND VPWR VPWR _13167_/X sky130_fd_sc_hd__mux2_2
X_10379_ _10379_/A VGND VGND VPWR VPWR _10379_/X sky130_fd_sc_hd__buf_1
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12118_ _12634_/A _12117_/A _12643_/A _12117_/Y VGND VGND VPWR VPWR _12640_/A sky130_fd_sc_hd__o22a_1
XFILLER_111_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13098_ _15644_/Q data_address[9] _15667_/Q VGND VGND VPWR VPWR _13098_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12049_ _12049_/A VGND VGND VPWR VPWR _12977_/A sky130_fd_sc_hd__buf_1
XFILLER_77_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07590_ _07591_/A _13075_/X VGND VGND VPWR VPWR _15490_/D sky130_fd_sc_hd__and2_1
XFILLER_37_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09260_ _15115_/Q _09249_/X _09259_/X _09252_/X VGND VGND VPWR VPWR _15115_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08211_ _08211_/A VGND VGND VPWR VPWR _08216_/A sky130_fd_sc_hd__clkbuf_2
X_09191_ _09199_/A VGND VGND VPWR VPWR _09191_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08142_ _08148_/A VGND VGND VPWR VPWR _08142_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08073_ _14309_/Q VGND VGND VPWR VPWR _08074_/A sky130_fd_sc_hd__buf_1
XFILLER_146_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08975_ _09007_/A VGND VGND VPWR VPWR _08994_/A sky130_fd_sc_hd__buf_2
XFILLER_29_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07926_ _07947_/A VGND VGND VPWR VPWR _07927_/A sky130_fd_sc_hd__buf_1
XFILLER_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07857_ _07786_/A _07709_/X _07871_/A _07774_/C _07710_/X VGND VGND VPWR VPWR _07863_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07788_ _07666_/Y _07668_/Y _07785_/Y _07787_/Y VGND VGND VPWR VPWR _07789_/B sky130_fd_sc_hd__a31o_1
XFILLER_83_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09527_ _10297_/A VGND VGND VPWR VPWR _09527_/X sky130_fd_sc_hd__buf_1
XFILLER_25_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ _09476_/A VGND VGND VPWR VPWR _09458_/X sky130_fd_sc_hd__buf_1
XFILLER_101_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08409_ _08409_/A VGND VGND VPWR VPWR _08409_/X sky130_fd_sc_hd__buf_1
XFILLER_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09389_ _09391_/A VGND VGND VPWR VPWR _09389_/X sky130_fd_sc_hd__clkbuf_1
X_11420_ _11422_/A VGND VGND VPWR VPWR _11420_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11351_ _11353_/A VGND VGND VPWR VPWR _11351_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10302_ _10302_/A VGND VGND VPWR VPWR _10302_/X sky130_fd_sc_hd__clkbuf_1
X_14070_ _14969_/Q _15065_/Q _15033_/Q _15097_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14070_/X sky130_fd_sc_hd__mux4_1
X_11282_ _11290_/A VGND VGND VPWR VPWR _11282_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13021_ _14365_/Q VGND VGND VPWR VPWR _13021_/Y sky130_fd_sc_hd__inv_2
X_10233_ _14869_/Q _10227_/X _09991_/X _10229_/X VGND VGND VPWR VPWR _14869_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10164_ _10164_/A VGND VGND VPWR VPWR _10171_/A sky130_fd_sc_hd__buf_1
XFILLER_105_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10095_ _10104_/A VGND VGND VPWR VPWR _10102_/A sky130_fd_sc_hd__buf_1
X_14972_ _09836_/X _14972_/D VGND VGND VPWR VPWR _14972_/Q sky130_fd_sc_hd__dfxtp_1
X_13923_ _14663_/Q _15239_/Q _14727_/Q _14695_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13923_/X sky130_fd_sc_hd__mux4_2
XFILLER_47_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13854_ _15182_/Q _15150_/Q _14766_/Q _14798_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13854_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12805_ _12805_/A VGND VGND VPWR VPWR _12805_/X sky130_fd_sc_hd__buf_1
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13785_ _15125_/Q _15349_/Q _15317_/Q _15285_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13785_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10997_ _11016_/A VGND VGND VPWR VPWR _10997_/X sky130_fd_sc_hd__buf_1
XFILLER_31_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15524_ _15527_/CLK _15524_/D VGND VGND VPWR VPWR _15524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12736_ _12736_/A _15573_/Q VGND VGND VPWR VPWR _12913_/A sky130_fd_sc_hd__nor2_2
XFILLER_31_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15455_ _15663_/CLK _15455_/D VGND VGND VPWR VPWR data_address[28] sky130_fd_sc_hd__dfxtp_4
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _12666_/X _12139_/X _12616_/X VGND VGND VPWR VPWR _12667_/Y sky130_fd_sc_hd__o21ai_2
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ _12008_/X _14406_/D VGND VGND VPWR VPWR _14406_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11618_ _14519_/Q _11612_/X _11484_/X _11613_/X VGND VGND VPWR VPWR _14519_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15386_ _08139_/X _15386_/D VGND VGND VPWR VPWR _15386_/Q sky130_fd_sc_hd__dfxtp_1
X_12598_ _12598_/A _12598_/B VGND VGND VPWR VPWR _12598_/Y sky130_fd_sc_hd__nor2_1
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14337_ _12018_/X _15671_/Q VGND VGND VPWR VPWR _14337_/Q sky130_fd_sc_hd__dfxtp_4
X_11549_ _11549_/A VGND VGND VPWR VPWR _11549_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14268_ _14501_/Q _14469_/Q _14437_/Q _14405_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14268_/X sky130_fd_sc_hd__mux4_2
XFILLER_143_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13219_ _13218_/X _12861_/X _15565_/Q VGND VGND VPWR VPWR _13219_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14199_ _14828_/Q _14860_/Q _14892_/Q _14924_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14199_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08760_ _15240_/Q _08753_/X _08517_/X _08754_/X VGND VGND VPWR VPWR _15240_/D sky130_fd_sc_hd__a22o_1
X_07711_ _13138_/X VGND VGND VPWR VPWR _07711_/X sky130_fd_sc_hd__buf_1
X_08691_ _15261_/Q _08679_/X _08384_/X _08682_/X VGND VGND VPWR VPWR _15261_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07642_ _07642_/A _15507_/Q VGND VGND VPWR VPWR _15459_/D sky130_fd_sc_hd__or2_1
XFILLER_38_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07573_ _07573_/A VGND VGND VPWR VPWR _07582_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09312_ _09312_/A VGND VGND VPWR VPWR _09376_/A sky130_fd_sc_hd__buf_2
XFILLER_34_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09243_ _09269_/A VGND VGND VPWR VPWR _09254_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09174_ _15135_/Q _09169_/X _09170_/X _09173_/X VGND VGND VPWR VPWR _15135_/D sky130_fd_sc_hd__a22o_1
X_08125_ _08144_/A VGND VGND VPWR VPWR _08125_/X sky130_fd_sc_hd__buf_1
XFILLER_147_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08056_ _08071_/A VGND VGND VPWR VPWR _08067_/A sky130_fd_sc_hd__buf_1
XFILLER_134_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08958_ _15195_/Q _08954_/X _08817_/X _08955_/X VGND VGND VPWR VPWR _15195_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07909_ _07908_/X _07909_/B _07909_/C VGND VGND VPWR VPWR _15428_/D sky130_fd_sc_hd__and3b_1
XFILLER_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08889_ _08894_/A VGND VGND VPWR VPWR _08889_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10920_ _10920_/A VGND VGND VPWR VPWR _10920_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10851_ _10851_/A VGND VGND VPWR VPWR _10913_/A sky130_fd_sc_hd__buf_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13570_ _13569_/X _14324_/D _15506_/Q VGND VGND VPWR VPWR _13570_/X sky130_fd_sc_hd__mux2_2
XFILLER_71_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10782_ _11528_/A VGND VGND VPWR VPWR _10782_/X sky130_fd_sc_hd__clkbuf_2
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12521_ _12860_/A _12521_/B VGND VGND VPWR VPWR _12521_/X sky130_fd_sc_hd__or2_1
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15240_ _08759_/X _15240_/D VGND VGND VPWR VPWR _15240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12452_ _12452_/A _12452_/B VGND VGND VPWR VPWR _12452_/X sky130_fd_sc_hd__or2_1
X_11403_ _11403_/A VGND VGND VPWR VPWR _11403_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15171_ _09036_/X _15171_/D VGND VGND VPWR VPWR _15171_/Q sky130_fd_sc_hd__dfxtp_1
X_12383_ _12451_/A VGND VGND VPWR VPWR _12383_/X sky130_fd_sc_hd__buf_1
XFILLER_153_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14122_ _15219_/Q _14547_/Q _14995_/Q _15411_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14122_/X sky130_fd_sc_hd__mux4_2
X_11334_ _11395_/A VGND VGND VPWR VPWR _11355_/A sky130_fd_sc_hd__buf_2
XFILLER_4_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14053_ _14682_/Q _15258_/Q _14746_/Q _14714_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14053_/X sky130_fd_sc_hd__mux4_2
XFILLER_113_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11265_ _11274_/A VGND VGND VPWR VPWR _11265_/X sky130_fd_sc_hd__buf_1
X_13004_ _14348_/Q VGND VGND VPWR VPWR _13004_/Y sky130_fd_sc_hd__inv_2
X_10216_ _10216_/A VGND VGND VPWR VPWR _10216_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11196_ _14629_/Q _11186_/X _11195_/X _11188_/X VGND VGND VPWR VPWR _14629_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10147_ _10166_/A VGND VGND VPWR VPWR _10147_/X sky130_fd_sc_hd__buf_1
XFILLER_48_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14955_ _09895_/X _14955_/D VGND VGND VPWR VPWR _14955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10078_ _10078_/A VGND VGND VPWR VPWR _10078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13906_ _13902_/X _13903_/X _13904_/X _13905_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13906_/X sky130_fd_sc_hd__mux4_2
X_14886_ _10169_/X _14886_/D VGND VGND VPWR VPWR _14886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13837_ _14640_/Q _14608_/Q _14576_/Q _15376_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13837_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13768_ _14519_/Q _14487_/Q _14455_/Q _14423_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13768_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15507_ _15604_/CLK _15507_/D VGND VGND VPWR VPWR _15507_/Q sky130_fd_sc_hd__dfxtp_1
X_12719_ _13244_/X _12707_/X _12711_/X _12717_/Y _12718_/Y VGND VGND VPWR VPWR _12719_/Y
+ sky130_fd_sc_hd__o2111ai_4
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_13699_ _14846_/Q _14878_/Q _14910_/Q _14942_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13699_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15438_ _15646_/CLK _15438_/D VGND VGND VPWR VPWR data_address[11] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15369_ _08198_/X _15369_/D VGND VGND VPWR VPWR _15369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09930_ _09945_/A VGND VGND VPWR VPWR _09931_/A sky130_fd_sc_hd__buf_1
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09861_ _09917_/A VGND VGND VPWR VPWR _09880_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08812_ _08825_/A VGND VGND VPWR VPWR _08812_/X sky130_fd_sc_hd__buf_1
XFILLER_140_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09792_ _09792_/A VGND VGND VPWR VPWR _09792_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08743_ _08743_/A VGND VGND VPWR VPWR _08763_/A sky130_fd_sc_hd__buf_1
XFILLER_39_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08674_ _08676_/A VGND VGND VPWR VPWR _08674_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07625_ _12035_/B VGND VGND VPWR VPWR _12984_/C sky130_fd_sc_hd__buf_1
XFILLER_42_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07556_ _07556_/A _07556_/B _07556_/C VGND VGND VPWR VPWR _12993_/A sky130_fd_sc_hd__and3_1
XFILLER_22_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07487_ _07573_/A VGND VGND VPWR VPWR _07569_/A sky130_fd_sc_hd__buf_1
XFILLER_139_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09226_ _15123_/Q _09223_/X _09224_/X _09225_/X VGND VGND VPWR VPWR _15123_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09157_ _15138_/Q _09152_/X _09153_/X _09156_/X VGND VGND VPWR VPWR _15138_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08108_ _08120_/A VGND VGND VPWR VPWR _08109_/A sky130_fd_sc_hd__clkbuf_2
X_09088_ _15158_/Q _09085_/X _08839_/X _09087_/X VGND VGND VPWR VPWR _15158_/D sky130_fd_sc_hd__a22o_1
X_08039_ _08071_/A VGND VGND VPWR VPWR _08052_/A sky130_fd_sc_hd__buf_2
XFILLER_89_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11050_ _11054_/A VGND VGND VPWR VPWR _11050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10001_ _14931_/Q _09998_/X _09999_/X _10000_/X VGND VGND VPWR VPWR _14931_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14740_ _10744_/X _14740_/D VGND VGND VPWR VPWR _14740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11952_ _14423_/Q _11946_/X _07994_/A _11947_/X VGND VGND VPWR VPWR _14423_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10903_ _10909_/A VGND VGND VPWR VPWR _10903_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14671_ _11019_/X _14671_/D VGND VGND VPWR VPWR _14671_/Q sky130_fd_sc_hd__dfxtp_1
X_11883_ _11889_/A VGND VGND VPWR VPWR _11883_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13622_ _13621_/X _14311_/D _15506_/Q VGND VGND VPWR VPWR _13622_/X sky130_fd_sc_hd__mux2_2
XFILLER_83_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10834_ _10834_/A VGND VGND VPWR VPWR _10901_/A sky130_fd_sc_hd__buf_1
Xrepeater13 _14402_/Q VGND VGND VPWR VPWR _13946_/S1 sky130_fd_sc_hd__clkbuf_16
XFILLER_60_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater24 _13919_/S0 VGND VGND VPWR VPWR _13918_/S0 sky130_fd_sc_hd__buf_12
Xrepeater35 _14397_/Q VGND VGND VPWR VPWR _14266_/S0 sky130_fd_sc_hd__clkbuf_16
X_13553_ _13552_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13553_/X sky130_fd_sc_hd__mux2_1
X_10765_ _10765_/A VGND VGND VPWR VPWR _11514_/A sky130_fd_sc_hd__buf_2
Xrepeater46 _14268_/S0 VGND VGND VPWR VPWR _14238_/S0 sky130_fd_sc_hd__buf_12
X_12504_ _12498_/X _12951_/B _12501_/X _12503_/X VGND VGND VPWR VPWR _12504_/Y sky130_fd_sc_hd__o22ai_4
X_13484_ _13483_/X _13072_/X _14336_/Q VGND VGND VPWR VPWR _13484_/X sky130_fd_sc_hd__mux2_1
X_10696_ _10706_/A VGND VGND VPWR VPWR _10696_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15223_ _08833_/X _15223_/D VGND VGND VPWR VPWR _15223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12435_ _12446_/B VGND VGND VPWR VPWR _12435_/X sky130_fd_sc_hd__buf_2
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15154_ _09101_/X _15154_/D VGND VGND VPWR VPWR _15154_/Q sky130_fd_sc_hd__dfxtp_1
X_12366_ _12362_/X _12395_/A _12365_/X _13190_/X _12493_/A VGND VGND VPWR VPWR _12366_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_126_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14105_ _15125_/Q _15349_/Q _15317_/Q _15285_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14105_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11317_ _11317_/A _11317_/B VGND VGND VPWR VPWR _11330_/A sky130_fd_sc_hd__or2_2
XFILLER_126_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15085_ _09373_/X _15085_/D VGND VGND VPWR VPWR _15085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12297_ _15553_/Q VGND VGND VPWR VPWR _12329_/A sky130_fd_sc_hd__inv_2
XFILLER_113_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14036_ _14032_/X _14033_/X _14034_/X _14035_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14036_/X sky130_fd_sc_hd__mux4_2
XFILLER_4_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11248_ _11559_/A VGND VGND VPWR VPWR _11439_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11179_ _14633_/Q _11173_/X _11178_/X _11175_/X VGND VGND VPWR VPWR _14633_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14938_ _09968_/X _14938_/D VGND VGND VPWR VPWR _14938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14869_ _10232_/X _14869_/D VGND VGND VPWR VPWR _14869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07410_ _07411_/A _13563_/X VGND VGND VPWR VPWR _15583_/D sky130_fd_sc_hd__and2_1
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08390_ _09184_/A VGND VGND VPWR VPWR _08390_/X sky130_fd_sc_hd__buf_1
XFILLER_23_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07341_ _07341_/A VGND VGND VPWR VPWR _07341_/X sky130_fd_sc_hd__buf_1
XFILLER_50_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07272_ _07273_/A _07272_/B VGND VGND VPWR VPWR _15620_/D sky130_fd_sc_hd__nor2_1
X_09011_ _15180_/Q _09006_/X _08883_/X _09008_/X VGND VGND VPWR VPWR _15180_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09913_ _09915_/A VGND VGND VPWR VPWR _09913_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09844_ _14970_/Q _09837_/X _09574_/X _09838_/X VGND VGND VPWR VPWR _14970_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09775_ _09783_/A VGND VGND VPWR VPWR _09775_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08726_ _08735_/A VGND VGND VPWR VPWR _08731_/A sky130_fd_sc_hd__buf_1
XFILLER_100_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08657_ _08659_/A VGND VGND VPWR VPWR _08657_/X sky130_fd_sc_hd__clkbuf_1
X_07608_ _07608_/A _13062_/X VGND VGND VPWR VPWR _15477_/D sky130_fd_sc_hd__and2_1
X_08588_ _08588_/A VGND VGND VPWR VPWR _08588_/X sky130_fd_sc_hd__buf_1
XFILLER_14_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07539_ _15468_/Q VGND VGND VPWR VPWR _07539_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10550_ _10550_/A VGND VGND VPWR VPWR _10550_/X sky130_fd_sc_hd__buf_1
XFILLER_139_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09209_ _09248_/A VGND VGND VPWR VPWR _09235_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10481_ _10481_/A VGND VGND VPWR VPWR _10490_/A sky130_fd_sc_hd__buf_1
X_12220_ _12220_/A VGND VGND VPWR VPWR _12220_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12151_ _15544_/Q _12151_/B VGND VGND VPWR VPWR _12151_/Y sky130_fd_sc_hd__nor2_2
XFILLER_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11102_ _11128_/A VGND VGND VPWR VPWR _11111_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12082_ _12102_/A VGND VGND VPWR VPWR _12082_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11033_ _14668_/Q _11025_/X _10788_/X _11027_/X VGND VGND VPWR VPWR _14668_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12984_ _12984_/A _12984_/B _12984_/C VGND VGND VPWR VPWR _12984_/X sky130_fd_sc_hd__and3_1
XFILLER_18_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14723_ _10830_/X _14723_/D VGND VGND VPWR VPWR _14723_/Q sky130_fd_sc_hd__dfxtp_1
X_11935_ _11941_/A VGND VGND VPWR VPWR _11935_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14654_ _11086_/X _14654_/D VGND VGND VPWR VPWR _14654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11866_ _11866_/A VGND VGND VPWR VPWR _11866_/X sky130_fd_sc_hd__buf_1
X_13605_ _13604_/X _07310_/Y _13649_/S VGND VGND VPWR VPWR _13605_/X sky130_fd_sc_hd__mux2_1
X_10817_ _10817_/A VGND VGND VPWR VPWR _10817_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14585_ _11353_/X _14585_/D VGND VGND VPWR VPWR _14585_/Q sky130_fd_sc_hd__dfxtp_1
X_11797_ _11805_/A VGND VGND VPWR VPWR _11797_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13536_ _14006_/X _14011_/X _14387_/Q VGND VGND VPWR VPWR _13536_/X sky130_fd_sc_hd__mux2_1
X_10748_ _10754_/A VGND VGND VPWR VPWR _10748_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13467_ _13786_/X _13791_/X _13521_/S VGND VGND VPWR VPWR _13467_/X sky130_fd_sc_hd__mux2_1
X_10679_ _10689_/A VGND VGND VPWR VPWR _10679_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15206_ _08908_/X _15206_/D VGND VGND VPWR VPWR _15206_/Q sky130_fd_sc_hd__dfxtp_1
X_12418_ _12414_/X _12415_/X _12416_/X _13180_/X _12417_/X VGND VGND VPWR VPWR _12418_/X
+ sky130_fd_sc_hd__o32a_1
X_13398_ _13400_/X _13399_/X _13415_/S VGND VGND VPWR VPWR _13398_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15137_ _09158_/X _15137_/D VGND VGND VPWR VPWR _15137_/Q sky130_fd_sc_hd__dfxtp_1
X_12349_ _12578_/A VGND VGND VPWR VPWR _12349_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15068_ _09435_/X _15068_/D VGND VGND VPWR VPWR _15068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14019_ _14846_/Q _14878_/Q _14910_/Q _14942_/Q _14060_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14019_/X sky130_fd_sc_hd__mux4_1
X_07890_ _13146_/X _07742_/Y _07889_/Y VGND VGND VPWR VPWR _07891_/B sky130_fd_sc_hd__o21ai_1
XFILLER_68_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09560_ _15037_/Q _09544_/X _09559_/X _09549_/X VGND VGND VPWR VPWR _15037_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08511_ _09267_/A VGND VGND VPWR VPWR _08511_/X sky130_fd_sc_hd__buf_1
X_09491_ _09495_/A VGND VGND VPWR VPWR _09491_/X sky130_fd_sc_hd__clkbuf_1
X_08442_ _09220_/A VGND VGND VPWR VPWR _08442_/X sky130_fd_sc_hd__buf_1
XFILLER_24_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ _15327_/Q _08366_/X _08369_/X _08372_/X VGND VGND VPWR VPWR _15327_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07324_ _07341_/A VGND VGND VPWR VPWR _07324_/X sky130_fd_sc_hd__buf_1
XFILLER_32_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07255_ _07256_/A _07255_/B VGND VGND VPWR VPWR _15632_/D sky130_fd_sc_hd__nor2_1
XFILLER_136_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07186_ rst VGND VGND VPWR VPWR _07247_/A sky130_fd_sc_hd__buf_1
XFILLER_118_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A VGND VGND VPWR VPWR _14397_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09827_ _09888_/A VGND VGND VPWR VPWR _09847_/A sky130_fd_sc_hd__buf_2
XFILLER_74_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09758_ _14995_/Q _09756_/X _09612_/X _09757_/X VGND VGND VPWR VPWR _14995_/D sky130_fd_sc_hd__a22o_1
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08709_ _15255_/Q _08702_/X _08420_/X _08703_/X VGND VGND VPWR VPWR _15255_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09689_ _09693_/A VGND VGND VPWR VPWR _09689_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11720_ _14490_/Q _11713_/X _11471_/X _11714_/X VGND VGND VPWR VPWR _14490_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11651_ _11651_/A VGND VGND VPWR VPWR _11673_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10602_ _10606_/A VGND VGND VPWR VPWR _10602_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ _15544_/CLK pc[31] VGND VGND VPWR VPWR _14370_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ _14530_/Q _11578_/X _11431_/X _11581_/X VGND VGND VPWR VPWR _14530_/D sky130_fd_sc_hd__a22o_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _13409_/X _13405_/X _13408_/S VGND VGND VPWR VPWR _13321_/X sky130_fd_sc_hd__mux2_1
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10533_ _10542_/A VGND VGND VPWR VPWR _10540_/A sky130_fd_sc_hd__buf_1
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13252_ _13253_/X _13265_/X _15562_/Q VGND VGND VPWR VPWR _13252_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10464_ _10470_/A VGND VGND VPWR VPWR _10464_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12203_ _12275_/A VGND VGND VPWR VPWR _12773_/A sky130_fd_sc_hd__buf_1
XFILLER_136_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13183_ _13186_/X _13206_/X _13408_/S VGND VGND VPWR VPWR _13183_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10395_ _10395_/A VGND VGND VPWR VPWR _10420_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12134_ _12661_/A _12133_/A _12132_/X _12133_/Y VGND VGND VPWR VPWR _12135_/A sky130_fd_sc_hd__o22a_1
XFILLER_123_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12065_ _15583_/Q VGND VGND VPWR VPWR _12065_/X sky130_fd_sc_hd__buf_1
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11016_ _11016_/A VGND VGND VPWR VPWR _11016_/X sky130_fd_sc_hd__buf_1
XFILLER_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12967_ _12967_/A _12967_/B VGND VGND VPWR VPWR _12967_/X sky130_fd_sc_hd__or2_1
XFILLER_33_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14706_ _10897_/X _14706_/D VGND VGND VPWR VPWR _14706_/Q sky130_fd_sc_hd__dfxtp_1
X_11918_ _14433_/Q _11912_/X _07936_/A _11915_/X VGND VGND VPWR VPWR _14433_/D sky130_fd_sc_hd__a22o_1
X_12898_ _12444_/Y _12447_/Y _12902_/C VGND VGND VPWR VPWR _12905_/B sky130_fd_sc_hd__o21bai_1
XFILLER_60_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11849_ _14453_/Q _11844_/X _08006_/A _11846_/X VGND VGND VPWR VPWR _14453_/D sky130_fd_sc_hd__a22o_1
X_14637_ _11158_/X _14637_/D VGND VGND VPWR VPWR _14637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14568_ _11411_/X _14568_/D VGND VGND VPWR VPWR _14568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13519_ _13518_/X rdata[1] _14338_/Q VGND VGND VPWR VPWR _13519_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14499_ _11683_/X _14499_/D VGND VGND VPWR VPWR _14499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08991_ _08991_/A VGND VGND VPWR VPWR _08998_/A sky130_fd_sc_hd__buf_1
XFILLER_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07942_ _07956_/A VGND VGND VPWR VPWR _07942_/X sky130_fd_sc_hd__buf_1
XFILLER_96_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07873_ _07873_/A VGND VGND VPWR VPWR _07878_/A sky130_fd_sc_hd__inv_2
XFILLER_110_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09612_ _10367_/A VGND VGND VPWR VPWR _09612_/X sky130_fd_sc_hd__buf_1
XFILLER_110_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09543_ _09640_/A VGND VGND VPWR VPWR _09577_/A sky130_fd_sc_hd__buf_2
XFILLER_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09474_ _09474_/A VGND VGND VPWR VPWR _09474_/X sky130_fd_sc_hd__clkbuf_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ _14323_/Q VGND VGND VPWR VPWR _10733_/A sky130_fd_sc_hd__buf_1
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _15329_/Q _08344_/X _08355_/X _08350_/X VGND VGND VPWR VPWR _15329_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07307_ _07307_/A VGND VGND VPWR VPWR _07373_/A sky130_fd_sc_hd__buf_1
X_08287_ _15346_/Q _08282_/X _08021_/X _08283_/X VGND VGND VPWR VPWR _15346_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07238_ _07240_/A _07246_/B _07242_/A _07286_/B VGND VGND VPWR VPWR _07239_/C sky130_fd_sc_hd__o31a_1
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07169_ _07265_/B _07169_/B VGND VGND VPWR VPWR _07205_/A sky130_fd_sc_hd__or2_1
XFILLER_106_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10180_ _10180_/A VGND VGND VPWR VPWR _10180_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13870_ _14957_/Q _15053_/Q _15021_/Q _15085_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13870_/X sky130_fd_sc_hd__mux4_2
XFILLER_47_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12821_ _12821_/A VGND VGND VPWR VPWR _12821_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15540_ _15544_/CLK _15540_/D VGND VGND VPWR VPWR _15540_/Q sky130_fd_sc_hd__dfxtp_1
X_12752_ _12752_/A VGND VGND VPWR VPWR _12752_/X sky130_fd_sc_hd__buf_1
XFILLER_15_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11703_ _11703_/A VGND VGND VPWR VPWR _11765_/A sky130_fd_sc_hd__buf_2
X_15471_ _15599_/CLK _15471_/D VGND VGND VPWR VPWR _15471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12683_ _13234_/X _12493_/X _12678_/X _12680_/X _12682_/X VGND VGND VPWR VPWR _12683_/Y
+ sky130_fd_sc_hd__o2111ai_4
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _11954_/X _14422_/D VGND VGND VPWR VPWR _14422_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11643_/A VGND VGND VPWR VPWR _11634_/X sky130_fd_sc_hd__buf_1
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14353_ _15621_/CLK pc[14] VGND VGND VPWR VPWR _14353_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _14533_/Q _11552_/X _11564_/X _11554_/X VGND VGND VPWR VPWR _14533_/D sky130_fd_sc_hd__a22o_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13304_ _12859_/Y _12797_/B _15563_/Q VGND VGND VPWR VPWR _13304_/X sky130_fd_sc_hd__mux2_1
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10516_ _10516_/A VGND VGND VPWR VPWR _10536_/A sky130_fd_sc_hd__clkbuf_2
X_14284_ _15171_/Q _15139_/Q _14755_/Q _14787_/Q _07387_/A _14284_/S1 VGND VGND VPWR
+ VPWR _14284_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11496_ _11508_/A VGND VGND VPWR VPWR _11505_/A sky130_fd_sc_hd__buf_1
XFILLER_109_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13235_ _13236_/X _13258_/X _13408_/S VGND VGND VPWR VPWR _13235_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10447_ _10447_/A VGND VGND VPWR VPWR _10447_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13166_ _13165_/X _13205_/X _13393_/S VGND VGND VPWR VPWR _13166_/X sky130_fd_sc_hd__mux2_1
X_10378_ _10378_/A VGND VGND VPWR VPWR _10378_/X sky130_fd_sc_hd__buf_1
X_12117_ _12117_/A VGND VGND VPWR VPWR _12117_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13097_ _15643_/Q data_address[8] _15667_/Q VGND VGND VPWR VPWR _13097_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12048_ _13425_/X VGND VGND VPWR VPWR _12048_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13999_ _14848_/Q _14880_/Q _14912_/Q _14944_/Q _07387_/A _14060_/S1 VGND VGND VPWR
+ VPWR _13999_/X sky130_fd_sc_hd__mux4_2
XFILLER_34_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15669_ _15669_/CLK _15669_/D VGND VGND VPWR VPWR _15669_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_190 _12812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08210_ _15365_/Q _08204_/X _08091_/X _08205_/X VGND VGND VPWR VPWR _15365_/D sky130_fd_sc_hd__a22o_1
X_09190_ _09190_/A VGND VGND VPWR VPWR _09199_/A sky130_fd_sc_hd__buf_1
XFILLER_119_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08141_ _08150_/A VGND VGND VPWR VPWR _08148_/A sky130_fd_sc_hd__buf_1
XFILLER_119_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08072_ _08082_/A VGND VGND VPWR VPWR _08072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08974_ _08993_/A VGND VGND VPWR VPWR _08974_/X sky130_fd_sc_hd__buf_1
XFILLER_114_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07925_ _09700_/A _11910_/A VGND VGND VPWR VPWR _07947_/A sky130_fd_sc_hd__or2_2
XFILLER_75_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07856_ _07856_/A VGND VGND VPWR VPWR _07871_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_83_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07787_ _07658_/A _07664_/X _07786_/X _13123_/X VGND VGND VPWR VPWR _07787_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09526_ _10664_/A VGND VGND VPWR VPWR _10297_/A sky130_fd_sc_hd__buf_1
XFILLER_71_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ _09487_/A VGND VGND VPWR VPWR _09476_/A sky130_fd_sc_hd__buf_2
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08408_ _09196_/A VGND VGND VPWR VPWR _08408_/X sky130_fd_sc_hd__buf_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09388_ _15082_/Q _09386_/X _09263_/X _09387_/X VGND VGND VPWR VPWR _15082_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08339_ _08352_/A VGND VGND VPWR VPWR _08339_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11350_ _14587_/Q _11343_/X _11099_/X _11344_/X VGND VGND VPWR VPWR _14587_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10301_ _14850_/Q _10296_/X _10297_/X _10300_/X VGND VGND VPWR VPWR _14850_/D sky130_fd_sc_hd__a22o_1
XFILLER_125_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11281_ _11301_/A VGND VGND VPWR VPWR _11290_/A sky130_fd_sc_hd__buf_1
XFILLER_106_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13020_ _14364_/Q VGND VGND VPWR VPWR _13020_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10232_ _10236_/A VGND VGND VPWR VPWR _10232_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10163_ _14888_/Q _10157_/X _10047_/X _10158_/X VGND VGND VPWR VPWR _14888_/D sky130_fd_sc_hd__a22o_1
XFILLER_120_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10094_ _14909_/Q _10086_/X _09954_/X _10089_/X VGND VGND VPWR VPWR _14909_/D sky130_fd_sc_hd__a22o_1
X_14971_ _09841_/X _14971_/D VGND VGND VPWR VPWR _14971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13922_ _15207_/Q _14535_/Q _14983_/Q _15399_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13922_/X sky130_fd_sc_hd__mux4_2
XFILLER_59_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13853_ _14670_/Q _15246_/Q _14734_/Q _14702_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13853_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12804_ _12264_/X _12803_/X _12264_/X _12803_/X VGND VGND VPWR VPWR _12804_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13784_ _15189_/Q _15157_/Q _14773_/Q _14805_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13784_/X sky130_fd_sc_hd__mux4_1
X_10996_ _11026_/A VGND VGND VPWR VPWR _11016_/A sky130_fd_sc_hd__buf_1
XFILLER_31_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15523_ _15527_/CLK _15523_/D VGND VGND VPWR VPWR _15523_/Q sky130_fd_sc_hd__dfxtp_1
X_12735_ _12735_/A _12735_/B VGND VGND VPWR VPWR _12735_/X sky130_fd_sc_hd__or2_1
XFILLER_16_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15454_ _15456_/CLK _15454_/D VGND VGND VPWR VPWR data_address[27] sky130_fd_sc_hd__dfxtp_4
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _15546_/Q VGND VGND VPWR VPWR _12666_/X sky130_fd_sc_hd__buf_1
XFILLER_31_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ _12010_/X _14405_/D VGND VGND VPWR VPWR _14405_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_opt_11_clk _14328_/CLK VGND VGND VPWR VPWR clkbuf_opt_11_clk/X sky130_fd_sc_hd__clkbuf_16
X_11617_ _11617_/A VGND VGND VPWR VPWR _11617_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _12578_/X _12587_/X _12589_/Y _12592_/X _12596_/X VGND VGND VPWR VPWR _12597_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_15385_ _08142_/X _15385_/D VGND VGND VPWR VPWR _15385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14336_ _12019_/X _15672_/Q VGND VGND VPWR VPWR _14336_/Q sky130_fd_sc_hd__dfxtp_4
X_11548_ _11556_/A VGND VGND VPWR VPWR _11548_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14267_ _14629_/Q _14597_/Q _14565_/Q _15365_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14267_/X sky130_fd_sc_hd__mux4_1
X_11479_ _11479_/A VGND VGND VPWR VPWR _11479_/X sky130_fd_sc_hd__buf_1
XFILLER_143_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13218_ _13220_/X _13263_/X _13393_/S VGND VGND VPWR VPWR _13218_/X sky130_fd_sc_hd__mux2_1
X_14198_ _14508_/Q _14476_/Q _14444_/Q _14412_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14198_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13149_ _12211_/X _12998_/Y _13152_/S VGND VGND VPWR VPWR _13149_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07710_ _07715_/A _13139_/X VGND VGND VPWR VPWR _07710_/X sky130_fd_sc_hd__or2_1
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08690_ _08692_/A VGND VGND VPWR VPWR _08690_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07641_ _07641_/A _15508_/Q VGND VGND VPWR VPWR _15460_/D sky130_fd_sc_hd__or2_1
XFILLER_38_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07572_ _07572_/A _13086_/X VGND VGND VPWR VPWR _15501_/D sky130_fd_sc_hd__and2_1
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09311_ _09335_/A VGND VGND VPWR VPWR _09311_/X sky130_fd_sc_hd__buf_1
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09242_ _09281_/A VGND VGND VPWR VPWR _09269_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09173_ _09197_/A VGND VGND VPWR VPWR _09173_/X sky130_fd_sc_hd__buf_1
XFILLER_119_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08124_ _08184_/A VGND VGND VPWR VPWR _08144_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_147_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08055_ _15404_/Q _08046_/X _08054_/X _08050_/X VGND VGND VPWR VPWR _15404_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08957_ _08959_/A VGND VGND VPWR VPWR _08957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07908_ _07910_/A _07760_/B _07760_/C VGND VGND VPWR VPWR _07908_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08888_ _15211_/Q _08877_/X _08887_/X _08880_/X VGND VGND VPWR VPWR _15211_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07839_ _07697_/A _07822_/A _07838_/X _07833_/A VGND VGND VPWR VPWR _15447_/D sky130_fd_sc_hd__o211a_1
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10850_ _10860_/A VGND VGND VPWR VPWR _10850_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09509_ _09603_/A VGND VGND VPWR VPWR _09536_/A sky130_fd_sc_hd__clkbuf_2
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10781_ _10781_/A VGND VGND VPWR VPWR _11528_/A sky130_fd_sc_hd__buf_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _12770_/A _12520_/B VGND VGND VPWR VPWR _12521_/B sky130_fd_sc_hd__or2_1
XFILLER_12_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _12451_/A VGND VGND VPWR VPWR _12451_/X sky130_fd_sc_hd__buf_1
XFILLER_138_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11402_ _14571_/Q _11394_/X _11170_/X _11396_/X VGND VGND VPWR VPWR _14571_/D sky130_fd_sc_hd__a22o_1
X_15170_ _09038_/X _15170_/D VGND VGND VPWR VPWR _15170_/Q sky130_fd_sc_hd__dfxtp_1
X_12382_ _12699_/B VGND VGND VPWR VPWR _12451_/A sky130_fd_sc_hd__buf_1
XANTENNA_90 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14121_ _14117_/X _14118_/X _14119_/X _14120_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14121_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11333_ _11333_/A VGND VGND VPWR VPWR _11395_/A sky130_fd_sc_hd__buf_2
XFILLER_126_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14052_ _15226_/Q _14554_/Q _15002_/Q _15418_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14052_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11264_ _11273_/A VGND VGND VPWR VPWR _11264_/X sky130_fd_sc_hd__buf_1
XFILLER_137_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13003_ _14347_/Q VGND VGND VPWR VPWR _13003_/Y sky130_fd_sc_hd__inv_2
X_10215_ _14874_/Q _10207_/X _09969_/X _10208_/X VGND VGND VPWR VPWR _14874_/D sky130_fd_sc_hd__a22o_1
X_11195_ _11564_/A VGND VGND VPWR VPWR _11195_/X sky130_fd_sc_hd__buf_1
XFILLER_67_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10146_ _10146_/A VGND VGND VPWR VPWR _10166_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10077_ _14913_/Q _10071_/X _09934_/X _10074_/X VGND VGND VPWR VPWR _14913_/D sky130_fd_sc_hd__a22o_1
X_14954_ _09897_/X _14954_/D VGND VGND VPWR VPWR _14954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13905_ _15113_/Q _15337_/Q _15305_/Q _15273_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13905_/X sky130_fd_sc_hd__mux4_1
X_14885_ _10171_/X _14885_/D VGND VGND VPWR VPWR _14885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13836_ _13832_/X _13833_/X _13834_/X _13835_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13836_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10979_ _10988_/A VGND VGND VPWR VPWR _10984_/A sky130_fd_sc_hd__buf_1
X_13767_ _14647_/Q _14615_/Q _14583_/Q _15383_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13767_/X sky130_fd_sc_hd__mux4_2
XFILLER_43_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15506_ _07934_/A _15506_/D VGND VGND VPWR VPWR _15506_/Q sky130_fd_sc_hd__dfxtp_4
X_12718_ _12689_/A _12689_/B _12512_/X _12690_/B VGND VGND VPWR VPWR _12718_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_149_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13698_ _14526_/Q _14494_/Q _14462_/Q _14430_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13698_/X sky130_fd_sc_hd__mux4_1
X_15437_ _15601_/CLK _15437_/D VGND VGND VPWR VPWR data_address[10] sky130_fd_sc_hd__dfxtp_4
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ _13328_/X _12620_/X _12593_/X _12648_/Y VGND VGND VPWR VPWR _12649_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15368_ _08200_/X _15368_/D VGND VGND VPWR VPWR _15368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14319_ _15599_/CLK _14319_/D VGND VGND VPWR VPWR _14319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15299_ _08542_/X _15299_/D VGND VGND VPWR VPWR _15299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09860_ _09860_/A VGND VGND VPWR VPWR _09917_/A sky130_fd_sc_hd__buf_2
XFILLER_97_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08811_ _08816_/A VGND VGND VPWR VPWR _08811_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09791_ _14985_/Q _09787_/X _09667_/X _09788_/X VGND VGND VPWR VPWR _14985_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08742_ _08762_/A VGND VGND VPWR VPWR _08742_/X sky130_fd_sc_hd__buf_1
XFILLER_85_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08673_ _15265_/Q _08666_/X _08355_/X _08669_/X VGND VGND VPWR VPWR _15265_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07624_ _15519_/Q VGND VGND VPWR VPWR _12035_/B sky130_fd_sc_hd__inv_2
XFILLER_26_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07555_ _07630_/B _07533_/A _07629_/B _14402_/Q _07554_/X VGND VGND VPWR VPWR _07556_/C
+ sky130_fd_sc_hd__o221a_1
X_07486_ _07486_/A _13517_/X VGND VGND VPWR VPWR _15531_/D sky130_fd_sc_hd__and2_1
XFILLER_139_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09225_ _09237_/A VGND VGND VPWR VPWR _09225_/X sky130_fd_sc_hd__buf_1
X_09156_ _09156_/A VGND VGND VPWR VPWR _09156_/X sky130_fd_sc_hd__buf_1
X_08107_ _09296_/A _11061_/A VGND VGND VPWR VPWR _08120_/A sky130_fd_sc_hd__or2_2
XFILLER_108_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09087_ _09107_/A VGND VGND VPWR VPWR _09087_/X sky130_fd_sc_hd__buf_1
XFILLER_108_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08038_ _08038_/A VGND VGND VPWR VPWR _08071_/A sky130_fd_sc_hd__buf_1
XFILLER_122_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10000_ _10013_/A VGND VGND VPWR VPWR _10000_/X sky130_fd_sc_hd__buf_1
X_09989_ _14934_/Q _09985_/X _09986_/X _09988_/X VGND VGND VPWR VPWR _14934_/D sky130_fd_sc_hd__a22o_1
XFILLER_76_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11951_ _11951_/A VGND VGND VPWR VPWR _11951_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10902_ _10922_/A VGND VGND VPWR VPWR _10909_/A sky130_fd_sc_hd__buf_1
X_11882_ _11900_/A VGND VGND VPWR VPWR _11889_/A sky130_fd_sc_hd__buf_1
X_14670_ _11021_/X _14670_/D VGND VGND VPWR VPWR _14670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13621_ _13620_/X _07343_/Y _13641_/S VGND VGND VPWR VPWR _13621_/X sky130_fd_sc_hd__mux2_1
X_10833_ _14723_/Q _10663_/A _10832_/X _10668_/A VGND VGND VPWR VPWR _14723_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater14 _14401_/Q VGND VGND VPWR VPWR _13966_/S0 sky130_fd_sc_hd__clkbuf_16
Xrepeater25 _13737_/S0 VGND VGND VPWR VPWR _13963_/S0 sky130_fd_sc_hd__clkbuf_16
X_10764_ _10764_/A VGND VGND VPWR VPWR _10764_/X sky130_fd_sc_hd__buf_1
Xrepeater36 _14060_/S1 VGND VGND VPWR VPWR _14057_/S1 sky130_fd_sc_hd__clkbuf_16
X_13552_ _14046_/X _14051_/X _14387_/Q VGND VGND VPWR VPWR _13552_/X sky130_fd_sc_hd__mux2_1
Xrepeater47 _14239_/S0 VGND VGND VPWR VPWR _14265_/S0 sky130_fd_sc_hd__buf_12
X_12503_ _12951_/A _12492_/X _12502_/X VGND VGND VPWR VPWR _12503_/X sky130_fd_sc_hd__o21a_1
X_13483_ _13482_/X rdata[13] _13516_/S VGND VGND VPWR VPWR _13483_/X sky130_fd_sc_hd__mux2_2
X_10695_ _10725_/A VGND VGND VPWR VPWR _10706_/A sky130_fd_sc_hd__buf_1
XFILLER_9_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12434_ _15557_/Q VGND VGND VPWR VPWR _12446_/B sky130_fd_sc_hd__inv_2
X_15222_ _08836_/X _15222_/D VGND VGND VPWR VPWR _15222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12365_ _12450_/A VGND VGND VPWR VPWR _12365_/X sky130_fd_sc_hd__clkbuf_2
X_15153_ _09103_/X _15153_/D VGND VGND VPWR VPWR _15153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14104_ _15189_/Q _15157_/Q _14773_/Q _14805_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14104_/X sky130_fd_sc_hd__mux4_1
X_11316_ _11316_/A VGND VGND VPWR VPWR _11316_/X sky130_fd_sc_hd__clkbuf_1
X_15084_ _09379_/X _15084_/D VGND VGND VPWR VPWR _15084_/Q sky130_fd_sc_hd__dfxtp_1
X_12296_ _12111_/Y _12144_/X _12637_/A _12295_/X VGND VGND VPWR VPWR _12432_/D sky130_fd_sc_hd__o31a_2
XFILLER_153_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14035_ _15132_/Q _15356_/Q _15324_/Q _15292_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14035_/X sky130_fd_sc_hd__mux4_2
XFILLER_107_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11247_ _14615_/Q _11241_/X _11116_/X _11242_/X VGND VGND VPWR VPWR _14615_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11178_ _11545_/A VGND VGND VPWR VPWR _11178_/X sky130_fd_sc_hd__buf_1
XFILLER_95_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10129_ _14899_/Q _10127_/X _09999_/X _10128_/X VGND VGND VPWR VPWR _14899_/D sky130_fd_sc_hd__a22o_1
X_14937_ _09971_/X _14937_/D VGND VGND VPWR VPWR _14937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14868_ _10234_/X _14868_/D VGND VGND VPWR VPWR _14868_/Q sky130_fd_sc_hd__dfxtp_1
X_13819_ _14834_/Q _14866_/Q _14898_/Q _14930_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13819_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14799_ _10508_/X _14799_/D VGND VGND VPWR VPWR _14799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07340_ _14390_/Q VGND VGND VPWR VPWR _07495_/B sky130_fd_sc_hd__inv_2
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07271_ _07273_/A _07271_/B VGND VGND VPWR VPWR _15621_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09010_ _09012_/A VGND VGND VPWR VPWR _09010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09912_ _14950_/Q _09907_/X _09682_/X _09908_/X VGND VGND VPWR VPWR _14950_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09843_ _09845_/A VGND VGND VPWR VPWR _09843_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09774_ _09785_/A VGND VGND VPWR VPWR _09783_/A sky130_fd_sc_hd__buf_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08725_ _15251_/Q _08723_/X _08448_/X _08724_/X VGND VGND VPWR VPWR _15251_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08656_ _15268_/Q _08552_/A _08540_/X _08555_/A VGND VGND VPWR VPWR _15268_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07607_ _07608_/A _13063_/X VGND VGND VPWR VPWR _15478_/D sky130_fd_sc_hd__and2_1
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08587_ _08587_/A VGND VGND VPWR VPWR _08587_/X sky130_fd_sc_hd__buf_1
X_07538_ _15468_/Q _07533_/Y _15470_/Q _07534_/Y _07537_/X VGND VGND VPWR VPWR _07545_/B
+ sky130_fd_sc_hd__o221a_1
X_07469_ _07469_/A VGND VGND VPWR VPWR _07472_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09208_ _09215_/A VGND VGND VPWR VPWR _09208_/X sky130_fd_sc_hd__clkbuf_1
X_10480_ _14807_/Q _10474_/X _10349_/X _10475_/X VGND VGND VPWR VPWR _14807_/D sky130_fd_sc_hd__a22o_1
X_09139_ _09146_/A VGND VGND VPWR VPWR _09144_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12150_ _12150_/A VGND VGND VPWR VPWR _12151_/B sky130_fd_sc_hd__inv_2
XFILLER_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11101_ _11101_/A VGND VGND VPWR VPWR _11128_/A sky130_fd_sc_hd__buf_1
X_12081_ _12081_/A VGND VGND VPWR VPWR _12102_/A sky130_fd_sc_hd__buf_1
XFILLER_151_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11032_ _11036_/A VGND VGND VPWR VPWR _11032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12983_ _15526_/Q _15527_/Q _12983_/C VGND VGND VPWR VPWR _12983_/Y sky130_fd_sc_hd__nor3_4
XFILLER_58_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14722_ _10837_/X _14722_/D VGND VGND VPWR VPWR _14722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11934_ _11934_/A VGND VGND VPWR VPWR _11941_/A sky130_fd_sc_hd__buf_1
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14653_ _11090_/X _14653_/D VGND VGND VPWR VPWR _14653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11865_ _11865_/A VGND VGND VPWR VPWR _11865_/X sky130_fd_sc_hd__buf_1
XFILLER_45_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13604_ _14176_/X _14181_/X _13648_/S VGND VGND VPWR VPWR _13604_/X sky130_fd_sc_hd__mux2_2
X_10816_ _14727_/Q _10812_/X _10814_/X _10815_/X VGND VGND VPWR VPWR _14727_/D sky130_fd_sc_hd__a22o_1
X_11796_ _14467_/Q _11688_/A _11570_/X _11691_/A VGND VGND VPWR VPWR _14467_/D sky130_fd_sc_hd__a22o_1
X_14584_ _11358_/X _14584_/D VGND VGND VPWR VPWR _14584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13535_ _13534_/X _13088_/X _14337_/Q VGND VGND VPWR VPWR _13535_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10747_ _14740_/Q _10732_/X _10746_/X _10736_/X VGND VGND VPWR VPWR _14740_/D sky130_fd_sc_hd__a22o_1
X_13466_ _13465_/X _13078_/X _14336_/Q VGND VGND VPWR VPWR _13466_/X sky130_fd_sc_hd__mux2_1
X_10678_ _14752_/Q _10663_/X _10677_/X _10668_/X VGND VGND VPWR VPWR _14752_/D sky130_fd_sc_hd__a22o_1
X_15205_ _08912_/X _15205_/D VGND VGND VPWR VPWR _15205_/Q sky130_fd_sc_hd__dfxtp_1
X_12417_ _12417_/A VGND VGND VPWR VPWR _12417_/X sky130_fd_sc_hd__buf_1
XFILLER_126_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13397_ _12435_/X _12480_/B _13418_/S VGND VGND VPWR VPWR _13397_/X sky130_fd_sc_hd__mux2_1
X_15136_ _09163_/X _15136_/D VGND VGND VPWR VPWR _15136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12348_ _12663_/A VGND VGND VPWR VPWR _12578_/A sky130_fd_sc_hd__buf_1
XFILLER_114_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12279_ _12754_/A _12183_/A _12209_/A _12277_/Y _12278_/Y VGND VGND VPWR VPWR _12279_/X
+ sky130_fd_sc_hd__o221a_1
X_15067_ _09440_/X _15067_/D VGND VGND VPWR VPWR _15067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14018_ _14526_/Q _14494_/Q _14462_/Q _14430_/Q _14060_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14018_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08510_ _10803_/A VGND VGND VPWR VPWR _09267_/A sky130_fd_sc_hd__buf_1
X_09490_ _09499_/A VGND VGND VPWR VPWR _09495_/A sky130_fd_sc_hd__buf_1
XFILLER_36_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08441_ _10745_/A VGND VGND VPWR VPWR _09220_/A sky130_fd_sc_hd__buf_1
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08372_ _08409_/A VGND VGND VPWR VPWR _08372_/X sky130_fd_sc_hd__buf_1
X_07323_ _07297_/A _07301_/A _07307_/A _07322_/X VGND VGND VPWR VPWR _07341_/A sky130_fd_sc_hd__o211a_1
X_07254_ _07256_/A _07254_/B VGND VGND VPWR VPWR _15633_/D sky130_fd_sc_hd__nor2_1
XFILLER_149_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07185_ _13120_/X _07180_/Y _07250_/B _07180_/A _07184_/X VGND VGND VPWR VPWR _15666_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_145_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09826_ _09826_/A VGND VGND VPWR VPWR _09888_/A sky130_fd_sc_hd__buf_2
XFILLER_47_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09757_ _09768_/A VGND VGND VPWR VPWR _09757_/X sky130_fd_sc_hd__buf_1
XFILLER_55_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08708_ _08710_/A VGND VGND VPWR VPWR _08708_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09688_ _15013_/Q _09675_/X _09687_/X _09678_/X VGND VGND VPWR VPWR _15013_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08639_ _15274_/Q _08637_/X _08505_/X _08638_/X VGND VGND VPWR VPWR _15274_/D sky130_fd_sc_hd__a22o_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11650_ _11658_/A VGND VGND VPWR VPWR _11650_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10601_ _10610_/A VGND VGND VPWR VPWR _10606_/A sky130_fd_sc_hd__buf_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11581_ _11581_/A VGND VGND VPWR VPWR _11581_/X sky130_fd_sc_hd__buf_1
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _13402_/X _13398_/X _13408_/S VGND VGND VPWR VPWR _13320_/X sky130_fd_sc_hd__mux2_1
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ _14792_/Q _10526_/X _10415_/X _10527_/X VGND VGND VPWR VPWR _14792_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13251_ _13252_/X _13276_/X _15563_/Q VGND VGND VPWR VPWR _13251_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10463_ _10481_/A VGND VGND VPWR VPWR _10470_/A sky130_fd_sc_hd__buf_1
XFILLER_6_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12202_ _15538_/Q VGND VGND VPWR VPWR _12275_/A sky130_fd_sc_hd__inv_2
XFILLER_109_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13182_ _12415_/X _12388_/X _15561_/Q VGND VGND VPWR VPWR _13182_/X sky130_fd_sc_hd__mux2_1
X_10394_ _10394_/A VGND VGND VPWR VPWR _10394_/X sky130_fd_sc_hd__buf_1
XFILLER_123_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12133_ _12133_/A VGND VGND VPWR VPWR _12133_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12064_ _15551_/Q VGND VGND VPWR VPWR _12577_/A sky130_fd_sc_hd__inv_2
XFILLER_104_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11015_ _11015_/A VGND VGND VPWR VPWR _11015_/X sky130_fd_sc_hd__buf_1
XFILLER_49_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12966_ _12518_/B _12955_/B _12616_/A _12965_/X VGND VGND VPWR VPWR _12966_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_45_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14705_ _10899_/X _14705_/D VGND VGND VPWR VPWR _14705_/Q sky130_fd_sc_hd__dfxtp_1
X_11917_ _11919_/A VGND VGND VPWR VPWR _11917_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12897_ _12463_/X _12470_/X _12473_/A _12466_/A VGND VGND VPWR VPWR _12902_/C sky130_fd_sc_hd__o22a_1
XFILLER_60_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14636_ _11165_/X _14636_/D VGND VGND VPWR VPWR _14636_/Q sky130_fd_sc_hd__dfxtp_1
X_11848_ _11848_/A VGND VGND VPWR VPWR _11848_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14567_ _11413_/X _14567_/D VGND VGND VPWR VPWR _14567_/Q sky130_fd_sc_hd__dfxtp_1
X_11779_ _14473_/Q _11774_/X _11545_/X _11775_/X VGND VGND VPWR VPWR _14473_/D sky130_fd_sc_hd__a22o_1
XFILLER_146_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13518_ _13956_/X _13961_/X _13521_/S VGND VGND VPWR VPWR _13518_/X sky130_fd_sc_hd__mux2_1
X_14498_ _11685_/X _14498_/D VGND VGND VPWR VPWR _14498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13449_ _13726_/X _13731_/X _14386_/Q VGND VGND VPWR VPWR _13449_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15119_ _09239_/X _15119_/D VGND VGND VPWR VPWR _15119_/Q sky130_fd_sc_hd__dfxtp_1
X_08990_ _15185_/Q _08984_/X _08861_/X _08985_/X VGND VGND VPWR VPWR _15185_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07941_ _07975_/A VGND VGND VPWR VPWR _07956_/A sky130_fd_sc_hd__buf_1
X_07872_ _07872_/A _07872_/B _07872_/C VGND VGND VPWR VPWR _15439_/D sky130_fd_sc_hd__and3_1
XFILLER_68_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09611_ _10750_/A VGND VGND VPWR VPWR _10367_/A sky130_fd_sc_hd__buf_1
XFILLER_28_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09542_ _09542_/A VGND VGND VPWR VPWR _09640_/A sky130_fd_sc_hd__buf_2
XFILLER_64_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09473_ _15057_/Q _09466_/X _09232_/X _09467_/X VGND VGND VPWR VPWR _15057_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08424_ _08463_/A VGND VGND VPWR VPWR _08424_/X sky130_fd_sc_hd__buf_1
XFILLER_24_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ _09159_/A VGND VGND VPWR VPWR _08355_/X sky130_fd_sc_hd__buf_1
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07306_ _14377_/Q _14376_/Q _07306_/C VGND VGND VPWR VPWR _07307_/A sky130_fd_sc_hd__or3_1
X_08286_ _08290_/A VGND VGND VPWR VPWR _08286_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07237_ _07237_/A VGND VGND VPWR VPWR _07246_/B sky130_fd_sc_hd__buf_1
XFILLER_153_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07168_ _07267_/B _07208_/A VGND VGND VPWR VPWR _07169_/B sky130_fd_sc_hd__or2_4
XFILLER_105_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09809_ _09809_/A VGND VGND VPWR VPWR _09809_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12820_ _12820_/A VGND VGND VPWR VPWR _12820_/X sky130_fd_sc_hd__buf_4
XFILLER_74_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12751_ _12193_/A _12750_/X _12193_/A _12750_/X VGND VGND VPWR VPWR _12751_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11702_ _11722_/A VGND VGND VPWR VPWR _11702_/X sky130_fd_sc_hd__buf_1
X_15470_ _15517_/CLK _15470_/D VGND VGND VPWR VPWR _15470_/Q sky130_fd_sc_hd__dfxtp_1
X_12682_ _12637_/Y _12135_/A _12581_/X _12144_/B _12681_/X VGND VGND VPWR VPWR _12682_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14421_ _11960_/X _14421_/D VGND VGND VPWR VPWR _14421_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11642_/A VGND VGND VPWR VPWR _11633_/X sky130_fd_sc_hd__buf_1
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14352_ _15667_/CLK pc[13] VGND VGND VPWR VPWR _14352_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ _11564_/A VGND VGND VPWR VPWR _11564_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _13351_/X _13349_/X _13408_/S VGND VGND VPWR VPWR _13303_/X sky130_fd_sc_hd__mux2_1
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10515_ _10535_/A VGND VGND VPWR VPWR _10515_/X sky130_fd_sc_hd__buf_1
XFILLER_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11495_ _14549_/Q _11488_/X _11494_/X _11491_/X VGND VGND VPWR VPWR _14549_/D sky130_fd_sc_hd__a22o_1
X_14283_ _14659_/Q _15235_/Q _14723_/Q _14691_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14283_/X sky130_fd_sc_hd__mux4_2
XFILLER_6_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13234_ _13233_/X _12967_/X _15565_/Q VGND VGND VPWR VPWR _13234_/X sky130_fd_sc_hd__mux2_2
X_10446_ _14817_/Q _10440_/X _10303_/X _10443_/X VGND VGND VPWR VPWR _14817_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10377_ _10382_/A VGND VGND VPWR VPWR _10377_/X sky130_fd_sc_hd__clkbuf_1
X_13165_ _13164_/X _13186_/X _13408_/S VGND VGND VPWR VPWR _13165_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12116_ _15548_/Q VGND VGND VPWR VPWR _12643_/A sky130_fd_sc_hd__buf_1
X_13096_ _15642_/Q data_address[7] _15667_/Q VGND VGND VPWR VPWR _13096_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12047_ _12324_/A VGND VGND VPWR VPWR _12316_/B sky130_fd_sc_hd__inv_2
XFILLER_77_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13998_ _14528_/Q _14496_/Q _14464_/Q _14432_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13998_/X sky130_fd_sc_hd__mux4_2
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12949_ _12949_/A _12949_/B VGND VGND VPWR VPWR _12949_/X sky130_fd_sc_hd__or2_1
XFILLER_33_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15668_ _15668_/CLK _15668_/D VGND VGND VPWR VPWR _15668_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_180 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 _12812_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR clkbuf_opt_8_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14619_ _11235_/X _14619_/D VGND VGND VPWR VPWR _14619_/Q sky130_fd_sc_hd__dfxtp_1
X_15599_ _15599_/CLK _15599_/D VGND VGND VPWR VPWR _15599_/Q sky130_fd_sc_hd__dfxtp_1
X_08140_ _15386_/Q _08134_/X _07978_/X _08135_/X VGND VGND VPWR VPWR _15386_/D sky130_fd_sc_hd__a22o_1
X_08071_ _08071_/A VGND VGND VPWR VPWR _08082_/A sky130_fd_sc_hd__buf_1
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08973_ _09005_/A VGND VGND VPWR VPWR _08993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07924_ _09922_/A VGND VGND VPWR VPWR _11910_/A sky130_fd_sc_hd__buf_1
XFILLER_84_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07855_ _07777_/D _07854_/Y _07838_/X _07849_/X VGND VGND VPWR VPWR _15443_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07786_ _07786_/A VGND VGND VPWR VPWR _07786_/X sky130_fd_sc_hd__buf_1
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09525_ _09525_/A VGND VGND VPWR VPWR _09525_/X sky130_fd_sc_hd__buf_1
XFILLER_36_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09456_ _09475_/A VGND VGND VPWR VPWR _09456_/X sky130_fd_sc_hd__buf_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08407_ _10717_/A VGND VGND VPWR VPWR _09196_/A sky130_fd_sc_hd__buf_1
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09387_ _09396_/A VGND VGND VPWR VPWR _09387_/X sky130_fd_sc_hd__buf_1
X_08338_ _15331_/Q _08227_/A _08099_/X _08230_/A VGND VGND VPWR VPWR _15331_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08269_ _15351_/Q _08261_/X _07994_/X _08262_/X VGND VGND VPWR VPWR _15351_/D sky130_fd_sc_hd__a22o_1
XFILLER_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10300_ _10300_/A VGND VGND VPWR VPWR _10300_/X sky130_fd_sc_hd__buf_1
XFILLER_137_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11280_ _11310_/A VGND VGND VPWR VPWR _11301_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10231_ _10231_/A VGND VGND VPWR VPWR _10236_/A sky130_fd_sc_hd__buf_2
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10162_ _10162_/A VGND VGND VPWR VPWR _10162_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10093_ _10093_/A VGND VGND VPWR VPWR _10093_/X sky130_fd_sc_hd__clkbuf_1
X_14970_ _09843_/X _14970_/D VGND VGND VPWR VPWR _14970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13921_ _13917_/X _13918_/X _13919_/X _13920_/X _14401_/Q _13966_/S1 VGND VGND VPWR
+ VPWR _13921_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13852_ _15214_/Q _14542_/Q _14990_/Q _15406_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13852_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12803_ _12803_/A _12803_/B VGND VGND VPWR VPWR _12803_/X sky130_fd_sc_hd__and2_1
XFILLER_74_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13783_ _14677_/Q _15253_/Q _14741_/Q _14709_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13783_/X sky130_fd_sc_hd__mux4_2
X_10995_ _11015_/A VGND VGND VPWR VPWR _10995_/X sky130_fd_sc_hd__buf_1
X_15522_ _15527_/CLK _15522_/D VGND VGND VPWR VPWR _15522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12734_ _13304_/X VGND VGND VPWR VPWR _12846_/A sky130_fd_sc_hd__inv_2
XFILLER_15_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15453_ _15663_/CLK _15453_/D VGND VGND VPWR VPWR data_address[26] sky130_fd_sc_hd__dfxtp_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12665_ _12636_/X _12664_/X _12636_/X _12664_/X VGND VGND VPWR VPWR _12665_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_70_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _12013_/X _14404_/D VGND VGND VPWR VPWR _14404_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _14520_/Q _11612_/X _11479_/X _11613_/X VGND VGND VPWR VPWR _14520_/D sky130_fd_sc_hd__a22o_1
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15384_ _08146_/X _15384_/D VGND VGND VPWR VPWR _15384_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12596_ _13292_/X _12368_/X _12593_/X _12595_/Y VGND VGND VPWR VPWR _12596_/X sky130_fd_sc_hd__o22a_1
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14335_ _15505_/CLK _14335_/D VGND VGND VPWR VPWR _14335_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11547_ _11547_/A VGND VGND VPWR VPWR _11556_/A sky130_fd_sc_hd__buf_1
XFILLER_144_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14266_ _14262_/X _14263_/X _14264_/X _14265_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14266_/X sky130_fd_sc_hd__mux4_2
X_11478_ _11478_/A VGND VGND VPWR VPWR _11478_/X sky130_fd_sc_hd__clkbuf_1
X_13217_ _12611_/X _12634_/X _13418_/S VGND VGND VPWR VPWR _13217_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10429_ _14821_/Q _10418_/X _10428_/X _10420_/X VGND VGND VPWR VPWR _14821_/D sky130_fd_sc_hd__a22o_1
X_14197_ _14636_/Q _14604_/Q _14572_/Q _15372_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14197_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13148_ _12838_/X _12999_/Y _13152_/S VGND VGND VPWR VPWR _13148_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13079_ _12633_/X _15581_/Q _13090_/S VGND VGND VPWR VPWR _13079_/X sky130_fd_sc_hd__mux2_1
X_07640_ _07640_/A _15509_/Q VGND VGND VPWR VPWR _15461_/D sky130_fd_sc_hd__and2_1
XFILLER_81_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07571_ _07572_/A _13087_/X VGND VGND VPWR VPWR _15502_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_45_clk _14315_/CLK VGND VGND VPWR VPWR _15604_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09310_ _09374_/A VGND VGND VPWR VPWR _09335_/A sky130_fd_sc_hd__buf_2
XFILLER_34_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09241_ _15119_/Q _09235_/X _09240_/X _09237_/X VGND VGND VPWR VPWR _15119_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09172_ _09251_/A VGND VGND VPWR VPWR _09197_/A sky130_fd_sc_hd__buf_2
X_08123_ _08123_/A VGND VGND VPWR VPWR _08184_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08054_ _08054_/A VGND VGND VPWR VPWR _08054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08956_ _15196_/Q _08954_/X _08813_/X _08955_/X VGND VGND VPWR VPWR _15196_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07907_ _13152_/X VGND VGND VPWR VPWR _07910_/A sky130_fd_sc_hd__buf_1
XFILLER_57_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08887_ _09259_/A VGND VGND VPWR VPWR _08887_/X sky130_fd_sc_hd__buf_1
XFILLER_84_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07838_ _07838_/A VGND VGND VPWR VPWR _07838_/X sky130_fd_sc_hd__buf_1
XFILLER_72_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07769_ _07769_/A _15600_/Q VGND VGND VPWR VPWR _07769_/X sky130_fd_sc_hd__or2_1
XFILLER_71_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_36_clk _14397_/CLK VGND VGND VPWR VPWR _15544_/CLK sky130_fd_sc_hd__clkbuf_16
X_09508_ _09508_/A VGND VGND VPWR VPWR _09603_/A sky130_fd_sc_hd__buf_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10780_ _10812_/A VGND VGND VPWR VPWR _10780_/X sky130_fd_sc_hd__buf_1
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09439_ _09439_/A VGND VGND VPWR VPWR _09444_/A sky130_fd_sc_hd__buf_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _12450_/A VGND VGND VPWR VPWR _12450_/X sky130_fd_sc_hd__buf_1
X_11401_ _11403_/A VGND VGND VPWR VPWR _11401_/X sky130_fd_sc_hd__clkbuf_1
X_12381_ _12904_/B VGND VGND VPWR VPWR _12381_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_80 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14120_ _14964_/Q _15060_/Q _15028_/Q _15092_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14120_/X sky130_fd_sc_hd__mux4_2
XFILLER_125_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11332_ _11354_/A VGND VGND VPWR VPWR _11332_/X sky130_fd_sc_hd__buf_1
XFILLER_153_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14051_ _14047_/X _14048_/X _14049_/X _14050_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14051_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11263_ _11269_/A VGND VGND VPWR VPWR _11263_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13002_ _14346_/Q VGND VGND VPWR VPWR _13002_/Y sky130_fd_sc_hd__inv_2
X_10214_ _10216_/A VGND VGND VPWR VPWR _10214_/X sky130_fd_sc_hd__clkbuf_1
X_11194_ _11200_/A VGND VGND VPWR VPWR _11194_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10145_ _10153_/A VGND VGND VPWR VPWR _10145_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10076_ _10078_/A VGND VGND VPWR VPWR _10076_/X sky130_fd_sc_hd__clkbuf_1
X_14953_ _09902_/X _14953_/D VGND VGND VPWR VPWR _14953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13904_ _15177_/Q _15145_/Q _14761_/Q _14793_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13904_/X sky130_fd_sc_hd__mux4_2
XFILLER_47_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14884_ _10176_/X _14884_/D VGND VGND VPWR VPWR _14884_/Q sky130_fd_sc_hd__dfxtp_1
X_13835_ _15120_/Q _15344_/Q _15312_/Q _15280_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13835_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clk _14397_/CLK VGND VGND VPWR VPWR _15654_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13766_ _13762_/X _13763_/X _13764_/X _13765_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13766_/X sky130_fd_sc_hd__mux4_2
X_10978_ _14684_/Q _10976_/X _10703_/X _10977_/X VGND VGND VPWR VPWR _14684_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15505_ _15505_/CLK _15505_/D VGND VGND VPWR VPWR wdata[31] sky130_fd_sc_hd__dfxtp_2
X_12717_ _12155_/X _12712_/X _12713_/X _12716_/X VGND VGND VPWR VPWR _12717_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13697_ _14654_/Q _14622_/Q _14590_/Q _15390_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13697_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15436_ _15667_/CLK _15436_/D VGND VGND VPWR VPWR data_address[9] sky130_fd_sc_hd__dfxtp_2
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ _12908_/A VGND VGND VPWR VPWR _12648_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15367_ _08203_/X _15367_/D VGND VGND VPWR VPWR _15367_/Q sky130_fd_sc_hd__dfxtp_1
X_12579_ _12579_/A VGND VGND VPWR VPWR _12579_/X sky130_fd_sc_hd__buf_1
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14318_ _15597_/CLK _14318_/D VGND VGND VPWR VPWR _14318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15298_ _08549_/X _15298_/D VGND VGND VPWR VPWR _15298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14249_ _14823_/Q _14855_/Q _14887_/Q _14919_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14249_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08810_ _15229_/Q _08798_/X _08809_/X _08802_/X VGND VGND VPWR VPWR _15229_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09790_ _09792_/A VGND VGND VPWR VPWR _09790_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08741_ _08741_/A VGND VGND VPWR VPWR _08762_/A sky130_fd_sc_hd__buf_1
XFILLER_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08672_ _08676_/A VGND VGND VPWR VPWR _08672_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07623_ _07626_/A _12980_/B VGND VGND VPWR VPWR _15472_/D sky130_fd_sc_hd__nor2_1
XFILLER_93_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk _14397_/CLK VGND VGND VPWR VPWR _15579_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07554_ _15515_/Q _07541_/Y _15514_/Q _07542_/Y VGND VGND VPWR VPWR _07554_/X sky130_fd_sc_hd__o22a_1
X_07485_ _07486_/A _13514_/X VGND VGND VPWR VPWR _15532_/D sky130_fd_sc_hd__and2_1
X_09224_ _09224_/A VGND VGND VPWR VPWR _09224_/X sky130_fd_sc_hd__buf_1
X_09155_ _09171_/A VGND VGND VPWR VPWR _09156_/A sky130_fd_sc_hd__buf_1
XFILLER_147_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08106_ _09923_/A _11574_/B _08925_/C VGND VGND VPWR VPWR _11061_/A sky130_fd_sc_hd__or3_1
XFILLER_147_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09086_ _09117_/A VGND VGND VPWR VPWR _09107_/A sky130_fd_sc_hd__clkbuf_2
X_08037_ _15407_/Q _08029_/X _08036_/X _08032_/X VGND VGND VPWR VPWR _15407_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09988_ _10013_/A VGND VGND VPWR VPWR _09988_/X sky130_fd_sc_hd__buf_1
XFILLER_107_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08939_ _08961_/A VGND VGND VPWR VPWR _08950_/A sky130_fd_sc_hd__buf_1
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11950_ _14424_/Q _11946_/X _07988_/A _11947_/X VGND VGND VPWR VPWR _14424_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10901_ _10901_/A VGND VGND VPWR VPWR _10922_/A sky130_fd_sc_hd__buf_4
XFILLER_84_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11881_ _11907_/A VGND VGND VPWR VPWR _11900_/A sky130_fd_sc_hd__buf_1
XFILLER_44_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13620_ _14216_/X _14221_/X _13648_/S VGND VGND VPWR VPWR _13620_/X sky130_fd_sc_hd__mux2_2
X_10832_ _11570_/A VGND VGND VPWR VPWR _10832_/X sky130_fd_sc_hd__buf_1
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater15 _14401_/Q VGND VGND VPWR VPWR _07533_/A sky130_fd_sc_hd__clkbuf_16
X_13551_ _13550_/X _13084_/X _14337_/Q VGND VGND VPWR VPWR _13551_/X sky130_fd_sc_hd__mux2_1
X_10763_ _10769_/A VGND VGND VPWR VPWR _10763_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater26 _13740_/S0 VGND VGND VPWR VPWR _13737_/S0 sky130_fd_sc_hd__clkbuf_16
Xrepeater37 _07379_/A VGND VGND VPWR VPWR _14060_/S1 sky130_fd_sc_hd__clkbuf_16
XFILLER_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater48 _14268_/S0 VGND VGND VPWR VPWR _14239_/S0 sky130_fd_sc_hd__clkbuf_16
X_12502_ _12714_/A VGND VGND VPWR VPWR _12502_/X sky130_fd_sc_hd__buf_1
XFILLER_40_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13482_ _13836_/X _13841_/X _13521_/S VGND VGND VPWR VPWR _13482_/X sky130_fd_sc_hd__mux2_2
XFILLER_139_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10694_ _10790_/A VGND VGND VPWR VPWR _10725_/A sky130_fd_sc_hd__buf_1
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15221_ _08843_/X _15221_/D VGND VGND VPWR VPWR _15221_/Q sky130_fd_sc_hd__dfxtp_1
X_12433_ _12415_/X _12407_/A _12429_/Y _12430_/Y _12432_/X VGND VGND VPWR VPWR _12443_/A
+ sky130_fd_sc_hd__o2111ai_4
X_15152_ _09105_/X _15152_/D VGND VGND VPWR VPWR _15152_/Q sky130_fd_sc_hd__dfxtp_1
X_12364_ _12478_/A VGND VGND VPWR VPWR _12450_/A sky130_fd_sc_hd__buf_1
XFILLER_4_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14103_ _14677_/Q _15253_/Q _14741_/Q _14709_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14103_/X sky130_fd_sc_hd__mux4_2
X_11315_ _14595_/Q _11207_/A _11201_/X _11210_/A VGND VGND VPWR VPWR _14595_/D sky130_fd_sc_hd__a22o_1
X_15083_ _09381_/X _15083_/D VGND VGND VPWR VPWR _15083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12295_ _12089_/Y _12286_/Y _12111_/Y _12292_/X _12294_/X VGND VGND VPWR VPWR _12295_/X
+ sky130_fd_sc_hd__o221a_1
X_14034_ _15196_/Q _15164_/Q _14780_/Q _14812_/Q _14055_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14034_/X sky130_fd_sc_hd__mux4_2
X_11246_ _11246_/A VGND VGND VPWR VPWR _11246_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11177_ _11177_/A VGND VGND VPWR VPWR _11177_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10128_ _10137_/A VGND VGND VPWR VPWR _10128_/X sky130_fd_sc_hd__buf_1
XFILLER_36_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10059_ _10428_/A VGND VGND VPWR VPWR _10059_/X sky130_fd_sc_hd__buf_1
X_14936_ _09976_/X _14936_/D VGND VGND VPWR VPWR _14936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14867_ _10236_/X _14867_/D VGND VGND VPWR VPWR _14867_/Q sky130_fd_sc_hd__dfxtp_1
X_13818_ _14514_/Q _14482_/Q _14450_/Q _14418_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13818_/X sky130_fd_sc_hd__mux4_2
XFILLER_23_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14798_ _10510_/X _14798_/D VGND VGND VPWR VPWR _14798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13749_ _14841_/Q _14873_/Q _14905_/Q _14937_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13749_/X sky130_fd_sc_hd__mux4_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07270_ _07270_/A VGND VGND VPWR VPWR _07273_/A sky130_fd_sc_hd__buf_1
X_15419_ _07971_/X _15419_/D VGND VGND VPWR VPWR _15419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_7_clk clkbuf_opt_5_clk/X VGND VGND VPWR VPWR _14391_/CLK sky130_fd_sc_hd__clkbuf_16
X_09911_ _09915_/A VGND VGND VPWR VPWR _09911_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09842_ _14971_/Q _09837_/X _09569_/X _09838_/X VGND VGND VPWR VPWR _14971_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09773_ _14990_/Q _09767_/X _09637_/X _09768_/X VGND VGND VPWR VPWR _14990_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08724_ _08733_/A VGND VGND VPWR VPWR _08724_/X sky130_fd_sc_hd__buf_1
XFILLER_85_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08655_ _08659_/A VGND VGND VPWR VPWR _08655_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07606_ _07608_/A _13064_/X VGND VGND VPWR VPWR _15479_/D sky130_fd_sc_hd__and2_1
XFILLER_82_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08586_ _08592_/A VGND VGND VPWR VPWR _08586_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07537_ _07535_/Y _07541_/A _15469_/Q _07536_/Y VGND VGND VPWR VPWR _07537_/X sky130_fd_sc_hd__o22a_1
X_07468_ _07468_/A _13481_/X VGND VGND VPWR VPWR _15543_/D sky130_fd_sc_hd__and2_1
XFILLER_50_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09207_ _15127_/Q _09195_/X _09206_/X _09197_/X VGND VGND VPWR VPWR _15127_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07399_ _07403_/A VGND VGND VPWR VPWR _07402_/A sky130_fd_sc_hd__clkbuf_1
X_09138_ _15143_/Q _09136_/X _08905_/X _09137_/X VGND VGND VPWR VPWR _15143_/D sky130_fd_sc_hd__a22o_1
X_09069_ _09089_/A VGND VGND VPWR VPWR _09074_/A sky130_fd_sc_hd__buf_1
X_11100_ _14651_/Q _11094_/X _11099_/X _11096_/X VGND VGND VPWR VPWR _14651_/D sky130_fd_sc_hd__a22o_1
XFILLER_150_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12080_ _12156_/A VGND VGND VPWR VPWR _12081_/A sky130_fd_sc_hd__buf_1
X_11031_ _11049_/A VGND VGND VPWR VPWR _11036_/A sky130_fd_sc_hd__buf_1
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12982_ _12982_/A VGND VGND VPWR VPWR _12982_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14721_ _10845_/X _14721_/D VGND VGND VPWR VPWR _14721_/Q sky130_fd_sc_hd__dfxtp_1
X_11933_ _14429_/Q _11925_/X _07963_/A _11928_/X VGND VGND VPWR VPWR _14429_/D sky130_fd_sc_hd__a22o_1
XFILLER_45_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14652_ _11093_/X _14652_/D VGND VGND VPWR VPWR _14652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11864_ _11868_/A VGND VGND VPWR VPWR _11864_/X sky130_fd_sc_hd__clkbuf_1
X_13603_ _13602_/X _13071_/X _14337_/Q VGND VGND VPWR VPWR _13603_/X sky130_fd_sc_hd__mux2_1
X_10815_ _10815_/A VGND VGND VPWR VPWR _10815_/X sky130_fd_sc_hd__buf_1
X_14583_ _11360_/X _14583_/D VGND VGND VPWR VPWR _14583_/Q sky130_fd_sc_hd__dfxtp_1
X_11795_ _11805_/A VGND VGND VPWR VPWR _11795_/X sky130_fd_sc_hd__clkbuf_1
X_13534_ _13533_/X _14333_/D _15506_/Q VGND VGND VPWR VPWR _13534_/X sky130_fd_sc_hd__mux2_1
X_10746_ _11498_/A VGND VGND VPWR VPWR _10746_/X sky130_fd_sc_hd__buf_1
XFILLER_41_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13465_ _13464_/X rdata[19] _13516_/S VGND VGND VPWR VPWR _13465_/X sky130_fd_sc_hd__mux2_2
X_10677_ _11443_/A VGND VGND VPWR VPWR _10677_/X sky130_fd_sc_hd__buf_1
XFILLER_139_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15204_ _08915_/X _15204_/D VGND VGND VPWR VPWR _15204_/Q sky130_fd_sc_hd__dfxtp_1
X_12416_ _12450_/A VGND VGND VPWR VPWR _12416_/X sky130_fd_sc_hd__buf_1
X_13396_ _12492_/X _12522_/X _15561_/Q VGND VGND VPWR VPWR _13396_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15135_ _09166_/X _15135_/D VGND VGND VPWR VPWR _15135_/Q sky130_fd_sc_hd__dfxtp_1
X_12347_ _12347_/A VGND VGND VPWR VPWR _12347_/X sky130_fd_sc_hd__buf_1
XFILLER_142_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15066_ _09442_/X _15066_/D VGND VGND VPWR VPWR _15066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12278_ _12752_/A _12183_/Y _12191_/Y VGND VGND VPWR VPWR _12278_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14017_ _14654_/Q _14622_/Q _14590_/Q _15390_/Q _14060_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14017_/X sky130_fd_sc_hd__mux4_2
X_11229_ _14621_/Q _11221_/X _11091_/X _11224_/X VGND VGND VPWR VPWR _14621_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14919_ _10049_/X _14919_/D VGND VGND VPWR VPWR _14919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08440_ _14321_/Q VGND VGND VPWR VPWR _10745_/A sky130_fd_sc_hd__buf_1
XFILLER_64_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08371_ _08486_/A VGND VGND VPWR VPWR _08409_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07322_ _07356_/A VGND VGND VPWR VPWR _07322_/X sky130_fd_sc_hd__buf_1
XFILLER_149_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07253_ _07257_/A VGND VGND VPWR VPWR _07256_/A sky130_fd_sc_hd__buf_1
X_07184_ _07184_/A VGND VGND VPWR VPWR _07184_/X sky130_fd_sc_hd__buf_1
XFILLER_129_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09825_ _09846_/A VGND VGND VPWR VPWR _09825_/X sky130_fd_sc_hd__buf_1
XFILLER_101_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09756_ _09767_/A VGND VGND VPWR VPWR _09756_/X sky130_fd_sc_hd__buf_1
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08707_ _15256_/Q _08702_/X _08414_/X _08703_/X VGND VGND VPWR VPWR _15256_/D sky130_fd_sc_hd__a22o_1
X_09687_ _10428_/A VGND VGND VPWR VPWR _09687_/X sky130_fd_sc_hd__buf_1
XFILLER_82_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08638_ _08648_/A VGND VGND VPWR VPWR _08638_/X sky130_fd_sc_hd__buf_1
XFILLER_82_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _15295_/Q _08565_/X _08369_/X _08568_/X VGND VGND VPWR VPWR _15295_/D sky130_fd_sc_hd__a22o_1
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ _14774_/Q _10597_/X _10354_/X _10599_/X VGND VGND VPWR VPWR _14774_/D sky130_fd_sc_hd__a22o_1
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11580_ _11592_/A VGND VGND VPWR VPWR _11581_/A sky130_fd_sc_hd__buf_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10531_ _10531_/A VGND VGND VPWR VPWR _10531_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13250_ _13251_/X _12846_/A _13393_/S VGND VGND VPWR VPWR _13250_/X sky130_fd_sc_hd__mux2_2
X_10462_ _10462_/A VGND VGND VPWR VPWR _10481_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_136_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12201_ _12201_/A VGND VGND VPWR VPWR _12209_/B sky130_fd_sc_hd__inv_2
X_13181_ _13182_/X _13192_/X _15562_/Q VGND VGND VPWR VPWR _13181_/X sky130_fd_sc_hd__mux2_1
X_10393_ _10418_/A VGND VGND VPWR VPWR _10393_/X sky130_fd_sc_hd__buf_1
XFILLER_109_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12132_ _15545_/Q VGND VGND VPWR VPWR _12132_/X sky130_fd_sc_hd__buf_1
XFILLER_108_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12063_ _12020_/X _12021_/X _12360_/A VGND VGND VPWR VPWR _12342_/A sky130_fd_sc_hd__o21a_1
XFILLER_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11014_ _11014_/A VGND VGND VPWR VPWR _11014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12965_ _12512_/A _12830_/A _12955_/Y VGND VGND VPWR VPWR _12965_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11916_ _14434_/Q _11912_/X _07929_/A _11915_/X VGND VGND VPWR VPWR _14434_/D sky130_fd_sc_hd__a22o_1
XFILLER_73_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14704_ _10903_/X _14704_/D VGND VGND VPWR VPWR _14704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12896_ _12951_/C _12896_/B VGND VGND VPWR VPWR _12905_/A sky130_fd_sc_hd__or2_2
XFILLER_61_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14635_ _11169_/X _14635_/D VGND VGND VPWR VPWR _14635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11847_ _14454_/Q _11844_/X _08000_/A _11846_/X VGND VGND VPWR VPWR _14454_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14566_ _11418_/X _14566_/D VGND VGND VPWR VPWR _14566_/Q sky130_fd_sc_hd__dfxtp_1
X_11778_ _11782_/A VGND VGND VPWR VPWR _11778_/X sky130_fd_sc_hd__clkbuf_1
X_13517_ _13516_/X _13061_/X _14336_/Q VGND VGND VPWR VPWR _13517_/X sky130_fd_sc_hd__mux2_1
X_10729_ _14743_/Q _10716_/X _10728_/X _10719_/X VGND VGND VPWR VPWR _14743_/D sky130_fd_sc_hd__a22o_1
X_14497_ _11695_/X _14497_/D VGND VGND VPWR VPWR _14497_/Q sky130_fd_sc_hd__dfxtp_1
X_13448_ _13447_/X _13084_/X _14336_/Q VGND VGND VPWR VPWR _13448_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13379_ _13381_/X _13380_/X _13415_/S VGND VGND VPWR VPWR _13379_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15118_ _09244_/X _15118_/D VGND VGND VPWR VPWR _15118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15049_ _09500_/X _15049_/D VGND VGND VPWR VPWR _15049_/Q sky130_fd_sc_hd__dfxtp_1
X_07940_ _08038_/A VGND VGND VPWR VPWR _07975_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07871_ _07871_/A _07871_/B VGND VGND VPWR VPWR _07872_/C sky130_fd_sc_hd__nand2_1
XFILLER_96_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09610_ _09625_/A VGND VGND VPWR VPWR _09610_/X sky130_fd_sc_hd__buf_1
XFILLER_95_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09541_ _09551_/A VGND VGND VPWR VPWR _09541_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09472_ _09474_/A VGND VGND VPWR VPWR _09472_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ _08481_/A VGND VGND VPWR VPWR _08463_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ _10671_/A VGND VGND VPWR VPWR _09159_/A sky130_fd_sc_hd__buf_1
X_07305_ _07306_/C VGND VGND VPWR VPWR _07321_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_149_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08285_ _08285_/A VGND VGND VPWR VPWR _08290_/A sky130_fd_sc_hd__buf_1
XFILLER_20_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07236_ _07236_/A VGND VGND VPWR VPWR _07240_/A sky130_fd_sc_hd__buf_1
X_07167_ _07268_/B _07167_/B VGND VGND VPWR VPWR _07208_/A sky130_fd_sc_hd__or2_1
XFILLER_3_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09808_ _14979_/Q _09702_/A _09695_/X _09705_/A VGND VGND VPWR VPWR _14979_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09739_ _09741_/A VGND VGND VPWR VPWR _09739_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12750_ _12750_/A _12750_/B VGND VGND VPWR VPWR _12750_/X sky130_fd_sc_hd__and2_1
XFILLER_55_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11701_ _11763_/A VGND VGND VPWR VPWR _11722_/A sky130_fd_sc_hd__buf_2
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12681_ _12681_/A VGND VGND VPWR VPWR _12681_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _11962_/X _14420_/D VGND VGND VPWR VPWR _14420_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11638_/A VGND VGND VPWR VPWR _11632_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14351_ _15647_/CLK pc[12] VGND VGND VPWR VPWR _14351_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ _11569_/A VGND VGND VPWR VPWR _11563_/X sky130_fd_sc_hd__buf_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _13348_/X _13346_/X _13408_/S VGND VGND VPWR VPWR _13302_/X sky130_fd_sc_hd__mux2_1
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10514_ _10514_/A VGND VGND VPWR VPWR _10535_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14282_ _15203_/Q _14531_/Q _14979_/Q _15395_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14282_/X sky130_fd_sc_hd__mux4_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11494_ _11494_/A VGND VGND VPWR VPWR _11494_/X sky130_fd_sc_hd__buf_1
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13233_ _13235_/X _13281_/X _13393_/S VGND VGND VPWR VPWR _13233_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10445_ _10447_/A VGND VGND VPWR VPWR _10445_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13164_ _13163_/X _13177_/X _13415_/S VGND VGND VPWR VPWR _13164_/X sky130_fd_sc_hd__mux2_1
X_10376_ _14833_/Q _10366_/X _10375_/X _10368_/X VGND VGND VPWR VPWR _14833_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12115_ _12113_/X _12103_/A _12645_/A _12084_/X VGND VGND VPWR VPWR _12117_/A sky130_fd_sc_hd__o22a_1
XFILLER_124_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13095_ _15641_/Q data_address[6] _15667_/Q VGND VGND VPWR VPWR _13095_/X sky130_fd_sc_hd__mux2_1
X_12046_ _12045_/Y _12031_/X _13424_/X _12024_/X _12041_/X VGND VGND VPWR VPWR _12324_/A
+ sky130_fd_sc_hd__o221a_2
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13997_ _14656_/Q _14624_/Q _14592_/Q _15392_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13997_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12948_ _12599_/X _12602_/X _12909_/A _12947_/X VGND VGND VPWR VPWR _12949_/B sky130_fd_sc_hd__o22a_1
XFILLER_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12879_ _12879_/A _12879_/B VGND VGND VPWR VPWR _12879_/Y sky130_fd_sc_hd__nand2_1
X_15667_ _15667_/CLK _15667_/D VGND VGND VPWR VPWR _15667_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_170 wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_181 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _12785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14618_ _11237_/X _14618_/D VGND VGND VPWR VPWR _14618_/Q sky130_fd_sc_hd__dfxtp_1
X_15598_ _15601_/CLK _15598_/D VGND VGND VPWR VPWR _15598_/Q sky130_fd_sc_hd__dfxtp_1
X_14549_ _11493_/X _14549_/D VGND VGND VPWR VPWR _14549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08070_ _15401_/Q _08062_/X _08069_/X _08065_/X VGND VGND VPWR VPWR _15401_/D sky130_fd_sc_hd__a22o_1
XFILLER_115_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08972_ _08980_/A VGND VGND VPWR VPWR _08972_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07923_ _08340_/B _08223_/B VGND VGND VPWR VPWR _09922_/A sky130_fd_sc_hd__or2_1
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07854_ _07854_/A VGND VGND VPWR VPWR _07854_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07785_ _07798_/A VGND VGND VPWR VPWR _07785_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09524_ _09542_/A VGND VGND VPWR VPWR _09525_/A sky130_fd_sc_hd__buf_1
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09455_ _09485_/A VGND VGND VPWR VPWR _09475_/A sky130_fd_sc_hd__buf_2
XFILLER_101_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08406_ _14326_/Q VGND VGND VPWR VPWR _10717_/A sky130_fd_sc_hd__buf_1
X_09386_ _09395_/A VGND VGND VPWR VPWR _09386_/X sky130_fd_sc_hd__buf_1
XFILLER_138_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08337_ _08352_/A VGND VGND VPWR VPWR _08337_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08268_ _08270_/A VGND VGND VPWR VPWR _08268_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07219_ _07273_/B _07163_/B _07212_/X _07217_/Y VGND VGND VPWR VPWR _15649_/D sky130_fd_sc_hd__a211oi_2
XFILLER_146_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08199_ _15369_/Q _08195_/X _08069_/X _08196_/X VGND VGND VPWR VPWR _15369_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10230_ _14870_/Q _10227_/X _09986_/X _10229_/X VGND VGND VPWR VPWR _14870_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10161_ _14889_/Q _10157_/X _10042_/X _10158_/X VGND VGND VPWR VPWR _14889_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10092_ _14910_/Q _10086_/X _09950_/X _10089_/X VGND VGND VPWR VPWR _14910_/D sky130_fd_sc_hd__a22o_1
XFILLER_120_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13920_ _14952_/Q _15048_/Q _15016_/Q _15080_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13920_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13851_ _13847_/X _13848_/X _13849_/X _13850_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13851_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12802_ _12802_/A _12802_/B VGND VGND VPWR VPWR _12803_/B sky130_fd_sc_hd__nand2_2
XFILLER_16_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13782_ _15221_/Q _14549_/Q _14997_/Q _15413_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13782_/X sky130_fd_sc_hd__mux4_1
X_10994_ _11024_/A VGND VGND VPWR VPWR _11015_/A sky130_fd_sc_hd__buf_1
XFILLER_16_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12733_ _13295_/X VGND VGND VPWR VPWR _12823_/A sky130_fd_sc_hd__inv_2
X_15521_ _15521_/CLK _15521_/D VGND VGND VPWR VPWR _15521_/Q sky130_fd_sc_hd__dfxtp_1
X_15452_ _15646_/CLK _15452_/D VGND VGND VPWR VPWR data_address[25] sky130_fd_sc_hd__dfxtp_2
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12662_/A _12133_/A _12581_/X _12144_/B VGND VGND VPWR VPWR _12664_/X sky130_fd_sc_hd__o22a_1
XFILLER_31_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _12015_/X _14403_/D VGND VGND VPWR VPWR _14403_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _11617_/A VGND VGND VPWR VPWR _11615_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15383_ _08148_/X _15383_/D VGND VGND VPWR VPWR _15383_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _12949_/A VGND VGND VPWR VPWR _12595_/Y sky130_fd_sc_hd__inv_2
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14334_ _15591_/CLK _14334_/D VGND VGND VPWR VPWR _14334_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ _14537_/Q _11540_/X _11545_/X _11542_/X VGND VGND VPWR VPWR _14537_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14265_ _15109_/Q _15333_/Q _15301_/Q _15269_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14265_/X sky130_fd_sc_hd__mux4_2
X_11477_ _14553_/Q _11474_/X _11475_/X _11476_/X VGND VGND VPWR VPWR _14553_/D sky130_fd_sc_hd__a22o_1
X_13216_ _13217_/X _13227_/X _13415_/S VGND VGND VPWR VPWR _13216_/X sky130_fd_sc_hd__mux2_1
X_10428_ _10428_/A VGND VGND VPWR VPWR _10428_/X sky130_fd_sc_hd__buf_1
X_14196_ _14192_/X _14193_/X _14194_/X _14195_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14196_/X sky130_fd_sc_hd__mux4_2
XFILLER_136_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13147_ _12847_/A _13000_/Y _13152_/S VGND VGND VPWR VPWR _13147_/X sky130_fd_sc_hd__mux2_1
X_10359_ _10359_/A VGND VGND VPWR VPWR _10359_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13078_ _12650_/Y _15580_/Q _13090_/S VGND VGND VPWR VPWR _13078_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12029_ _12050_/B VGND VGND VPWR VPWR _12029_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07570_ _07572_/A _13088_/X VGND VGND VPWR VPWR _15503_/D sky130_fd_sc_hd__and2_1
XFILLER_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09240_ _09240_/A VGND VGND VPWR VPWR _09240_/X sky130_fd_sc_hd__buf_1
X_09171_ _09171_/A VGND VGND VPWR VPWR _09251_/A sky130_fd_sc_hd__buf_2
X_08122_ _08143_/A VGND VGND VPWR VPWR _08122_/X sky130_fd_sc_hd__buf_1
X_08053_ _14313_/Q VGND VGND VPWR VPWR _08054_/A sky130_fd_sc_hd__buf_1
XFILLER_135_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08955_ _08964_/A VGND VGND VPWR VPWR _08955_/X sky130_fd_sc_hd__buf_1
XFILLER_88_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07906_ _07762_/A _07905_/A _07762_/Y _07905_/Y _07835_/X VGND VGND VPWR VPWR _15429_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08886_ _08894_/A VGND VGND VPWR VPWR _08886_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07837_ _07695_/Y _07833_/Y _07834_/Y _07835_/X _07836_/Y VGND VGND VPWR VPWR _15448_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_45_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07768_ _07897_/A _07752_/Y _07765_/Y _07767_/X VGND VGND VPWR VPWR _07889_/A sky130_fd_sc_hd__a31o_1
XFILLER_72_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09507_ _15047_/Q _09505_/X _09275_/X _09506_/X VGND VGND VPWR VPWR _15047_/D sky130_fd_sc_hd__a22o_1
X_07699_ _07832_/A _07834_/A VGND VGND VPWR VPWR _07778_/C sky130_fd_sc_hd__or2_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09438_ _15068_/Q _09436_/X _09184_/X _09437_/X VGND VGND VPWR VPWR _15068_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09369_ _15087_/Q _09365_/X _09240_/X _09366_/X VGND VGND VPWR VPWR _15087_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11400_ _14572_/Q _11394_/X _11166_/X _11396_/X VGND VGND VPWR VPWR _14572_/D sky130_fd_sc_hd__a22o_1
X_12380_ _12379_/A _12379_/B _12379_/Y VGND VGND VPWR VPWR _12904_/B sky130_fd_sc_hd__a21oi_2
XANTENNA_70 pc[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_81 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_92 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11331_ _11393_/A VGND VGND VPWR VPWR _11354_/A sky130_fd_sc_hd__buf_2
XFILLER_4_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14050_ _14971_/Q _15067_/Q _15035_/Q _15099_/Q _14395_/Q _14060_/S1 VGND VGND VPWR
+ VPWR _14050_/X sky130_fd_sc_hd__mux4_1
X_11262_ _11271_/A VGND VGND VPWR VPWR _11269_/A sky130_fd_sc_hd__buf_1
XFILLER_118_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13001_ _14345_/Q VGND VGND VPWR VPWR _13001_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10213_ _14875_/Q _10207_/X _09962_/X _10208_/X VGND VGND VPWR VPWR _14875_/D sky130_fd_sc_hd__a22o_1
X_11193_ _11203_/A VGND VGND VPWR VPWR _11200_/A sky130_fd_sc_hd__buf_1
XFILLER_106_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10144_ _10164_/A VGND VGND VPWR VPWR _10153_/A sky130_fd_sc_hd__buf_1
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A VGND VGND VPWR VPWR _14315_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10075_ _14914_/Q _10071_/X _09928_/X _10074_/X VGND VGND VPWR VPWR _14914_/D sky130_fd_sc_hd__a22o_1
X_14952_ _09904_/X _14952_/D VGND VGND VPWR VPWR _14952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13903_ _14665_/Q _15241_/Q _14729_/Q _14697_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13903_/X sky130_fd_sc_hd__mux4_2
XFILLER_36_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14883_ _10178_/X _14883_/D VGND VGND VPWR VPWR _14883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13834_ _15184_/Q _15152_/Q _14768_/Q _14800_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13834_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13765_ _15127_/Q _15351_/Q _15319_/Q _15287_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13765_/X sky130_fd_sc_hd__mux4_2
X_10977_ _10986_/A VGND VGND VPWR VPWR _10977_/X sky130_fd_sc_hd__buf_1
X_15504_ _15592_/CLK _15504_/D VGND VGND VPWR VPWR wdata[30] sky130_fd_sc_hd__dfxtp_2
XFILLER_149_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12716_ _12708_/X _12709_/X _12715_/X VGND VGND VPWR VPWR _12716_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13696_ _13692_/X _13693_/X _13694_/X _13695_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13696_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15435_ _15667_/CLK _15435_/D VGND VGND VPWR VPWR data_address[8] sky130_fd_sc_hd__dfxtp_4
X_12647_ _12643_/X _12113_/X _12634_/X _12645_/X VGND VGND VPWR VPWR _12908_/A sky130_fd_sc_hd__o22a_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15366_ _08207_/X _15366_/D VGND VGND VPWR VPWR _15366_/Q sky130_fd_sc_hd__dfxtp_1
X_12578_ _12578_/A VGND VGND VPWR VPWR _12578_/X sky130_fd_sc_hd__clkbuf_4
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14317_ _15668_/CLK _14317_/D VGND VGND VPWR VPWR _14317_/Q sky130_fd_sc_hd__dfxtp_1
X_11529_ _11529_/A VGND VGND VPWR VPWR _11554_/A sky130_fd_sc_hd__buf_1
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15297_ _08557_/X _15297_/D VGND VGND VPWR VPWR _15297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14248_ _14503_/Q _14471_/Q _14439_/Q _14407_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14248_/X sky130_fd_sc_hd__mux4_2
X_14179_ _14830_/Q _14862_/Q _14894_/Q _14926_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14179_/X sky130_fd_sc_hd__mux4_2
XFILLER_124_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08740_ _08740_/A VGND VGND VPWR VPWR _08740_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08671_ _08671_/A VGND VGND VPWR VPWR _08676_/A sky130_fd_sc_hd__buf_2
XFILLER_66_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07622_ _07622_/A VGND VGND VPWR VPWR _12980_/B sky130_fd_sc_hd__buf_1
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07553_ _15517_/Q VGND VGND VPWR VPWR _07629_/B sky130_fd_sc_hd__inv_2
XFILLER_81_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07484_ _07486_/A _13511_/X VGND VGND VPWR VPWR _15533_/D sky130_fd_sc_hd__and2_1
X_09223_ _09235_/A VGND VGND VPWR VPWR _09223_/X sky130_fd_sc_hd__buf_1
XFILLER_10_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09154_ _09167_/A VGND VGND VPWR VPWR _09171_/A sky130_fd_sc_hd__inv_2
XFILLER_148_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08105_ _11574_/A VGND VGND VPWR VPWR _09923_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_147_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09085_ _09106_/A VGND VGND VPWR VPWR _09085_/X sky130_fd_sc_hd__buf_1
X_08036_ _08036_/A VGND VGND VPWR VPWR _08036_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09987_ _10026_/A VGND VGND VPWR VPWR _10013_/A sky130_fd_sc_hd__buf_2
XFILLER_107_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08938_ _08970_/A VGND VGND VPWR VPWR _08961_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08869_ _09240_/A VGND VGND VPWR VPWR _08869_/X sky130_fd_sc_hd__buf_1
XFILLER_45_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10900_ _14705_/Q _10894_/X _10761_/X _10895_/X VGND VGND VPWR VPWR _14705_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11880_ _14444_/Q _11875_/X _08054_/A _11877_/X VGND VGND VPWR VPWR _14444_/D sky130_fd_sc_hd__a22o_1
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10831_ _10831_/A VGND VGND VPWR VPWR _11570_/A sky130_fd_sc_hd__buf_1
XFILLER_72_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13550_ _13549_/X _14329_/D _15506_/Q VGND VGND VPWR VPWR _13550_/X sky130_fd_sc_hd__mux2_1
X_10762_ _14737_/Q _10749_/X _10761_/X _10752_/X VGND VGND VPWR VPWR _14737_/D sky130_fd_sc_hd__a22o_1
Xrepeater16 _13950_/S1 VGND VGND VPWR VPWR _13860_/S1 sky130_fd_sc_hd__clkbuf_16
Xrepeater27 _07542_/A VGND VGND VPWR VPWR _13740_/S0 sky130_fd_sc_hd__clkbuf_16
XFILLER_40_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater38 _07379_/A VGND VGND VPWR VPWR _14284_/S1 sky130_fd_sc_hd__clkbuf_16
XFILLER_13_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12501_ _12753_/A VGND VGND VPWR VPWR _12501_/X sky130_fd_sc_hd__buf_2
XFILLER_13_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater49 _07387_/A VGND VGND VPWR VPWR _14268_/S0 sky130_fd_sc_hd__clkbuf_16
X_13481_ _13480_/X _13073_/X _14336_/Q VGND VGND VPWR VPWR _13481_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10693_ _10834_/A VGND VGND VPWR VPWR _10790_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_139_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15220_ _08847_/X _15220_/D VGND VGND VPWR VPWR _15220_/Q sky130_fd_sc_hd__dfxtp_1
X_12432_ _12432_/A _12432_/B _12432_/C _12432_/D VGND VGND VPWR VPWR _12432_/X sky130_fd_sc_hd__or4_4
XFILLER_12_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15151_ _09110_/X _15151_/D VGND VGND VPWR VPWR _15151_/Q sky130_fd_sc_hd__dfxtp_1
X_12363_ _12363_/A VGND VGND VPWR VPWR _12395_/A sky130_fd_sc_hd__buf_4
XFILLER_153_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14102_ _15221_/Q _14549_/Q _14997_/Q _15413_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14102_/X sky130_fd_sc_hd__mux4_1
X_11314_ _11316_/A VGND VGND VPWR VPWR _11314_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15082_ _09385_/X _15082_/D VGND VGND VPWR VPWR _15082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12294_ _12590_/A _12086_/A _12076_/A _12087_/Y VGND VGND VPWR VPWR _12294_/X sky130_fd_sc_hd__o22a_1
X_14033_ _14684_/Q _15260_/Q _14748_/Q _14716_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14033_/X sky130_fd_sc_hd__mux4_1
X_11245_ _14616_/Q _11241_/X _11112_/X _11242_/X VGND VGND VPWR VPWR _14616_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11176_ _14634_/Q _11173_/X _11174_/X _11175_/X VGND VGND VPWR VPWR _14634_/D sky130_fd_sc_hd__a22o_1
XFILLER_122_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10127_ _10136_/A VGND VGND VPWR VPWR _10127_/X sky130_fd_sc_hd__buf_1
XFILLER_67_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10058_ _10064_/A VGND VGND VPWR VPWR _10058_/X sky130_fd_sc_hd__clkbuf_1
X_14935_ _09980_/X _14935_/D VGND VGND VPWR VPWR _14935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14866_ _10242_/X _14866_/D VGND VGND VPWR VPWR _14866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13817_ _14642_/Q _14610_/Q _14578_/Q _15378_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13817_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14797_ _10513_/X _14797_/D VGND VGND VPWR VPWR _14797_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_opt_0_clk _14315_/CLK VGND VGND VPWR VPWR _14372_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13748_ _14521_/Q _14489_/Q _14457_/Q _14425_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13748_/X sky130_fd_sc_hd__mux4_2
XFILLER_149_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13679_ _14848_/Q _14880_/Q _14912_/Q _14944_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13679_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15418_ _07976_/X _15418_/D VGND VGND VPWR VPWR _15418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15349_ _08277_/X _15349_/D VGND VGND VPWR VPWR _15349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09910_ _09910_/A VGND VGND VPWR VPWR _09915_/A sky130_fd_sc_hd__buf_1
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09841_ _09845_/A VGND VGND VPWR VPWR _09841_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09772_ _09772_/A VGND VGND VPWR VPWR _09772_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08723_ _08732_/A VGND VGND VPWR VPWR _08723_/X sky130_fd_sc_hd__buf_1
X_08654_ _08671_/A VGND VGND VPWR VPWR _08659_/A sky130_fd_sc_hd__buf_1
X_07605_ _07609_/A VGND VGND VPWR VPWR _07608_/A sky130_fd_sc_hd__clkbuf_1
X_08585_ _08605_/A VGND VGND VPWR VPWR _08592_/A sky130_fd_sc_hd__buf_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07536_ _14402_/Q VGND VGND VPWR VPWR _07536_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07467_ _07468_/A _13478_/X VGND VGND VPWR VPWR _15544_/D sky130_fd_sc_hd__and2_1
X_09206_ _09206_/A VGND VGND VPWR VPWR _09206_/X sky130_fd_sc_hd__buf_1
XFILLER_22_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07398_ _07612_/A _13531_/X VGND VGND VPWR VPWR _15591_/D sky130_fd_sc_hd__and2_1
X_09137_ _09137_/A VGND VGND VPWR VPWR _09137_/X sky130_fd_sc_hd__buf_1
XFILLER_136_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09068_ _09068_/A VGND VGND VPWR VPWR _09089_/A sky130_fd_sc_hd__buf_2
XFILLER_118_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08019_ _08019_/A VGND VGND VPWR VPWR _08019_/X sky130_fd_sc_hd__clkbuf_1
X_11030_ _11101_/A VGND VGND VPWR VPWR _11049_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12981_ _07619_/B _12973_/C _12980_/X VGND VGND VPWR VPWR _12981_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14720_ _10847_/X _14720_/D VGND VGND VPWR VPWR _14720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11932_ _11932_/A VGND VGND VPWR VPWR _11932_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11863_ _14449_/Q _11856_/X _08026_/A _11857_/X VGND VGND VPWR VPWR _14449_/D sky130_fd_sc_hd__a22o_1
X_14651_ _11098_/X _14651_/D VGND VGND VPWR VPWR _14651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10814_ _11553_/A VGND VGND VPWR VPWR _10814_/X sky130_fd_sc_hd__buf_1
X_13602_ _13601_/X _14316_/D _15506_/Q VGND VGND VPWR VPWR _13602_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11794_ _11807_/A VGND VGND VPWR VPWR _11805_/A sky130_fd_sc_hd__buf_1
X_14582_ _11362_/X _14582_/D VGND VGND VPWR VPWR _14582_/Q sky130_fd_sc_hd__dfxtp_1
X_10745_ _10745_/A VGND VGND VPWR VPWR _11498_/A sky130_fd_sc_hd__clkbuf_2
X_13533_ _13532_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13533_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13464_ _13776_/X _13781_/X _13521_/S VGND VGND VPWR VPWR _13464_/X sky130_fd_sc_hd__mux2_1
X_10676_ _10676_/A VGND VGND VPWR VPWR _11443_/A sky130_fd_sc_hd__buf_1
XFILLER_9_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12415_ _12415_/A VGND VGND VPWR VPWR _12415_/X sky130_fd_sc_hd__buf_4
X_15203_ _08918_/X _15203_/D VGND VGND VPWR VPWR _15203_/Q sky130_fd_sc_hd__dfxtp_1
X_13395_ _13397_/X _13396_/X _13415_/S VGND VGND VPWR VPWR _13395_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12346_ _12346_/A VGND VGND VPWR VPWR _12347_/A sky130_fd_sc_hd__buf_1
X_15134_ _09175_/X _15134_/D VGND VGND VPWR VPWR _15134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15065_ _09444_/X _15065_/D VGND VGND VPWR VPWR _15065_/Q sky130_fd_sc_hd__dfxtp_1
X_12277_ _12277_/A VGND VGND VPWR VPWR _12277_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14016_ _14012_/X _14013_/X _14014_/X _14015_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14016_/X sky130_fd_sc_hd__mux4_2
X_11228_ _11228_/A VGND VGND VPWR VPWR _11228_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11159_ _11159_/A VGND VGND VPWR VPWR _11186_/A sky130_fd_sc_hd__buf_1
XFILLER_122_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14918_ _10054_/X _14918_/D VGND VGND VPWR VPWR _14918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14849_ _10302_/X _14849_/D VGND VGND VPWR VPWR _14849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08370_ _08370_/A VGND VGND VPWR VPWR _08486_/A sky130_fd_sc_hd__buf_4
XFILLER_51_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07321_ _07559_/C _07321_/B _07321_/C VGND VGND VPWR VPWR _07356_/A sky130_fd_sc_hd__or3_1
XFILLER_149_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07252_ _07252_/A _07252_/B VGND VGND VPWR VPWR _15634_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07183_ _07221_/A VGND VGND VPWR VPWR _07184_/A sky130_fd_sc_hd__buf_1
XFILLER_145_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09824_ _09886_/A VGND VGND VPWR VPWR _09846_/A sky130_fd_sc_hd__buf_2
XFILLER_140_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09755_ _09761_/A VGND VGND VPWR VPWR _09755_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08706_ _08710_/A VGND VGND VPWR VPWR _08706_/X sky130_fd_sc_hd__clkbuf_1
X_09686_ _10823_/A VGND VGND VPWR VPWR _10428_/A sky130_fd_sc_hd__buf_1
XFILLER_27_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08637_ _08647_/A VGND VGND VPWR VPWR _08637_/X sky130_fd_sc_hd__buf_1
XFILLER_82_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08568_ _08588_/A VGND VGND VPWR VPWR _08568_/X sky130_fd_sc_hd__buf_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07519_ _07568_/A _14373_/Q VGND VGND VPWR VPWR _15509_/D sky130_fd_sc_hd__and2_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ _09259_/A VGND VGND VPWR VPWR _08499_/X sky130_fd_sc_hd__buf_1
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10530_ _14793_/Q _10526_/X _10411_/X _10527_/X VGND VGND VPWR VPWR _14793_/D sky130_fd_sc_hd__a22o_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10461_ _14813_/Q _10453_/X _10324_/X _10456_/X VGND VGND VPWR VPWR _14813_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12200_ _12774_/A _12199_/A _12791_/A _12199_/Y VGND VGND VPWR VPWR _12201_/A sky130_fd_sc_hd__o22a_1
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13180_ _13179_/X _13262_/X _15565_/Q VGND VGND VPWR VPWR _13180_/X sky130_fd_sc_hd__mux2_1
X_10392_ _10392_/A VGND VGND VPWR VPWR _10418_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12131_ _15577_/Q _12092_/A _12675_/A _12130_/X VGND VGND VPWR VPWR _12133_/A sky130_fd_sc_hd__o22a_1
XFILLER_123_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12062_ _12500_/A VGND VGND VPWR VPWR _12360_/A sky130_fd_sc_hd__buf_1
XFILLER_150_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11013_ _14673_/Q _11006_/X _10761_/X _11007_/X VGND VGND VPWR VPWR _14673_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12964_ _12962_/Y _12952_/Y _12963_/X VGND VGND VPWR VPWR _12972_/A sky130_fd_sc_hd__o21ai_4
XFILLER_92_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14703_ _10907_/X _14703_/D VGND VGND VPWR VPWR _14703_/Q sky130_fd_sc_hd__dfxtp_1
X_11915_ _11915_/A VGND VGND VPWR VPWR _11915_/X sky130_fd_sc_hd__buf_1
X_12895_ _12498_/X _15559_/Q _12495_/A _12491_/A VGND VGND VPWR VPWR _12896_/B sky130_fd_sc_hd__o22a_1
XFILLER_33_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14634_ _11172_/X _14634_/D VGND VGND VPWR VPWR _14634_/Q sky130_fd_sc_hd__dfxtp_1
X_11846_ _11866_/A VGND VGND VPWR VPWR _11846_/X sky130_fd_sc_hd__buf_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11777_ _11777_/A VGND VGND VPWR VPWR _11782_/A sky130_fd_sc_hd__buf_1
X_14565_ _11420_/X _14565_/D VGND VGND VPWR VPWR _14565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10728_ _11484_/A VGND VGND VPWR VPWR _10728_/X sky130_fd_sc_hd__buf_1
X_13516_ _13515_/X rdata[2] _13516_/S VGND VGND VPWR VPWR _13516_/X sky130_fd_sc_hd__mux2_2
XFILLER_13_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14496_ _11697_/X _14496_/D VGND VGND VPWR VPWR _14496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13447_ _13446_/X rdata[25] _13516_/S VGND VGND VPWR VPWR _13447_/X sky130_fd_sc_hd__mux2_1
X_10659_ _14755_/Q _10550_/A _10434_/X _10553_/A VGND VGND VPWR VPWR _14755_/D sky130_fd_sc_hd__a22o_1
XFILLER_127_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13378_ _12730_/A _12709_/X _13418_/S VGND VGND VPWR VPWR _13378_/X sky130_fd_sc_hd__mux2_1
X_15117_ _09247_/X _15117_/D VGND VGND VPWR VPWR _15117_/Q sky130_fd_sc_hd__dfxtp_1
X_12329_ _12329_/A VGND VGND VPWR VPWR _12329_/X sky130_fd_sc_hd__buf_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15048_ _09502_/X _15048_/D VGND VGND VPWR VPWR _15048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07870_ _07868_/A _07867_/Y _07868_/Y _07867_/A _07869_/X VGND VGND VPWR VPWR _15440_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09540_ _15040_/Q _09525_/X _09539_/X _09530_/X VGND VGND VPWR VPWR _15040_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09471_ _15058_/Q _09466_/X _09228_/X _09467_/X VGND VGND VPWR VPWR _15058_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08422_ _08431_/A VGND VGND VPWR VPWR _08422_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08353_ _14334_/Q VGND VGND VPWR VPWR _10671_/A sky130_fd_sc_hd__buf_1
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07304_ _14375_/Q _07559_/B VGND VGND VPWR VPWR _07306_/C sky130_fd_sc_hd__or2_1
X_08284_ _15347_/Q _08282_/X _08016_/X _08283_/X VGND VGND VPWR VPWR _15347_/D sky130_fd_sc_hd__a22o_1
XFILLER_137_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07235_ _07235_/A VGND VGND VPWR VPWR _07288_/A sky130_fd_sc_hd__buf_1
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07166_ _07269_/B _07214_/A VGND VGND VPWR VPWR _07167_/B sky130_fd_sc_hd__or2_2
XFILLER_117_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09807_ _09809_/A VGND VGND VPWR VPWR _09807_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07999_ _14323_/Q VGND VGND VPWR VPWR _08000_/A sky130_fd_sc_hd__buf_1
XFILLER_101_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09738_ _15001_/Q _09736_/X _09579_/X _09737_/X VGND VGND VPWR VPWR _15001_/D sky130_fd_sc_hd__a22o_1
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09669_ _09684_/A VGND VGND VPWR VPWR _09680_/A sky130_fd_sc_hd__buf_1
XFILLER_70_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11700_ _11700_/A VGND VGND VPWR VPWR _11763_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12680_ _12662_/X _12676_/X _12384_/X _12679_/Y VGND VGND VPWR VPWR _12680_/X sky130_fd_sc_hd__a22o_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11649_/A VGND VGND VPWR VPWR _11638_/A sky130_fd_sc_hd__buf_1
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14350_ _15652_/CLK pc[11] VGND VGND VPWR VPWR _14350_/Q sky130_fd_sc_hd__dfxtp_1
X_11562_ _11587_/A VGND VGND VPWR VPWR _11569_/A sky130_fd_sc_hd__buf_1
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13301_ _13302_/X _12489_/B _13393_/S VGND VGND VPWR VPWR _13301_/X sky130_fd_sc_hd__mux2_2
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10513_ _10521_/A VGND VGND VPWR VPWR _10513_/X sky130_fd_sc_hd__clkbuf_1
X_14281_ _14277_/X _14278_/X _14279_/X _14280_/X _14397_/Q _14398_/Q VGND VGND VPWR
+ VPWR _14281_/X sky130_fd_sc_hd__mux4_1
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11493_ _11493_/A VGND VGND VPWR VPWR _11493_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13232_ _12138_/X _12662_/X _15561_/Q VGND VGND VPWR VPWR _13232_/X sky130_fd_sc_hd__mux2_1
X_10444_ _14818_/Q _10440_/X _10297_/X _10443_/X VGND VGND VPWR VPWR _14818_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13163_ _12492_/X _12480_/B _13418_/S VGND VGND VPWR VPWR _13163_/X sky130_fd_sc_hd__mux2_1
X_10375_ _10375_/A VGND VGND VPWR VPWR _10375_/X sky130_fd_sc_hd__buf_1
XFILLER_124_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12114_ _15580_/Q VGND VGND VPWR VPWR _12645_/A sky130_fd_sc_hd__inv_2
XFILLER_97_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13094_ _15640_/Q data_address[5] _15667_/Q VGND VGND VPWR VPWR _13094_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12045_ _13423_/X VGND VGND VPWR VPWR _12045_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13996_ _13992_/X _13993_/X _13994_/X _13995_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _13996_/X sky130_fd_sc_hd__mux4_2
X_12947_ _12615_/X _12618_/X _12909_/C _12945_/X _12946_/X VGND VGND VPWR VPWR _12947_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15666_ _15666_/CLK _15666_/D VGND VGND VPWR VPWR _15666_/Q sky130_fd_sc_hd__dfxtp_1
X_12878_ _12878_/A _12878_/B VGND VGND VPWR VPWR _12878_/X sky130_fd_sc_hd__or2_1
XANTENNA_160 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_182 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_193 _12480_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14617_ _11240_/X _14617_/D VGND VGND VPWR VPWR _14617_/Q sky130_fd_sc_hd__dfxtp_1
X_11829_ _14459_/Q _11825_/X _07973_/A _11826_/X VGND VGND VPWR VPWR _14459_/D sky130_fd_sc_hd__a22o_1
X_15597_ _15597_/CLK _15597_/D VGND VGND VPWR VPWR _15597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14548_ _11497_/X _14548_/D VGND VGND VPWR VPWR _14548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14479_ _11758_/X _14479_/D VGND VGND VPWR VPWR _14479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08971_ _08991_/A VGND VGND VPWR VPWR _08980_/A sky130_fd_sc_hd__buf_1
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07922_ _08778_/C _14299_/Q VGND VGND VPWR VPWR _08223_/B sky130_fd_sc_hd__or2b_1
XFILLER_69_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07853_ _07852_/A _07851_/Y _07852_/Y _07851_/A _07844_/X VGND VGND VPWR VPWR _15444_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07784_ _07803_/A _07808_/A _07804_/A _07804_/B _07783_/X VGND VGND VPWR VPWR _07798_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09523_ _10548_/A _09523_/B VGND VGND VPWR VPWR _09542_/A sky130_fd_sc_hd__or2_1
XFILLER_25_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09454_ _09454_/A VGND VGND VPWR VPWR _09454_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08405_ _08405_/A VGND VGND VPWR VPWR _08405_/X sky130_fd_sc_hd__buf_1
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09385_ _09391_/A VGND VGND VPWR VPWR _09385_/X sky130_fd_sc_hd__clkbuf_1
X_08336_ _08357_/A VGND VGND VPWR VPWR _08352_/A sky130_fd_sc_hd__buf_1
X_08267_ _15352_/Q _08261_/X _07988_/X _08262_/X VGND VGND VPWR VPWR _15352_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07218_ _13104_/X _07217_/Y _07209_/X _07165_/B VGND VGND VPWR VPWR _15650_/D sky130_fd_sc_hd__o211a_1
XFILLER_152_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08198_ _08200_/A VGND VGND VPWR VPWR _08198_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07149_ _13095_/X VGND VGND VPWR VPWR _07285_/B sky130_fd_sc_hd__inv_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10160_ _10162_/A VGND VGND VPWR VPWR _10160_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10091_ _10093_/A VGND VGND VPWR VPWR _10091_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13850_ _14959_/Q _15055_/Q _15023_/Q _15087_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13850_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12801_ _12798_/X _12839_/B _12839_/A _12267_/X VGND VGND VPWR VPWR _12802_/B sky130_fd_sc_hd__a31o_1
X_10993_ _10993_/A VGND VGND VPWR VPWR _10993_/X sky130_fd_sc_hd__buf_2
X_13781_ _13777_/X _13778_/X _13779_/X _13780_/X _07533_/A _14402_/Q VGND VGND VPWR
+ VPWR _13781_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15520_ _15521_/CLK _15520_/D VGND VGND VPWR VPWR _15520_/Q sky130_fd_sc_hd__dfxtp_1
X_12732_ _12460_/X _12723_/Y _12729_/Y _12731_/X VGND VGND VPWR VPWR _12732_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15451_ _15663_/CLK _15451_/D VGND VGND VPWR VPWR data_address[24] sky130_fd_sc_hd__dfxtp_1
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12663_ _12663_/A VGND VGND VPWR VPWR _12663_/X sky130_fd_sc_hd__buf_2
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14402_ _15648_/CLK instruction[18] VGND VGND VPWR VPWR _14402_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _14521_/Q _11612_/X _11475_/X _11613_/X VGND VGND VPWR VPWR _14521_/D sky130_fd_sc_hd__a22o_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ _08151_/X _15382_/D VGND VGND VPWR VPWR _15382_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _12588_/X _12079_/X _12590_/X _12591_/X VGND VGND VPWR VPWR _12949_/A sky130_fd_sc_hd__o22a_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14333_ _15498_/CLK _14333_/D VGND VGND VPWR VPWR _14333_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11545_ _11545_/A VGND VGND VPWR VPWR _11545_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14264_ _15173_/Q _15141_/Q _14757_/Q _14789_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14264_/X sky130_fd_sc_hd__mux4_1
X_11476_ _11476_/A VGND VGND VPWR VPWR _11476_/X sky130_fd_sc_hd__buf_1
XFILLER_109_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13215_ _13216_/X _13236_/X _13408_/S VGND VGND VPWR VPWR _13215_/X sky130_fd_sc_hd__mux2_1
X_10427_ _10433_/A VGND VGND VPWR VPWR _10427_/X sky130_fd_sc_hd__clkbuf_1
X_14195_ _15116_/Q _15340_/Q _15308_/Q _15276_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14195_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13146_ _12820_/X _13001_/Y _13152_/S VGND VGND VPWR VPWR _13146_/X sky130_fd_sc_hd__mux2_2
X_10358_ _10358_/A VGND VGND VPWR VPWR _10358_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13077_ _12660_/Y _15579_/Q _13090_/S VGND VGND VPWR VPWR _13077_/X sky130_fd_sc_hd__mux2_1
X_10289_ _14852_/Q _10183_/A _10062_/X _10186_/A VGND VGND VPWR VPWR _14852_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12028_ _07622_/A _15519_/Q _07617_/A _12974_/B VGND VGND VPWR VPWR _12050_/B sky130_fd_sc_hd__a31o_1
XFILLER_66_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13979_ _14850_/Q _14882_/Q _14914_/Q _14946_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _13979_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15649_ _15652_/CLK _15649_/D VGND VGND VPWR VPWR _15649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09170_ _09170_/A VGND VGND VPWR VPWR _09170_/X sky130_fd_sc_hd__buf_1
XFILLER_147_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08121_ _08182_/A VGND VGND VPWR VPWR _08143_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08052_ _08052_/A VGND VGND VPWR VPWR _08052_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08954_ _08963_/A VGND VGND VPWR VPWR _08954_/X sky130_fd_sc_hd__buf_1
XFILLER_57_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07905_ _07905_/A VGND VGND VPWR VPWR _07905_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08885_ _08885_/A VGND VGND VPWR VPWR _08894_/A sky130_fd_sc_hd__buf_1
X_07836_ _07695_/Y _07833_/Y _07834_/Y VGND VGND VPWR VPWR _07836_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07767_ _07746_/A _15598_/Q _07766_/X VGND VGND VPWR VPWR _07767_/X sky130_fd_sc_hd__a21bo_1
XFILLER_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09506_ _09506_/A VGND VGND VPWR VPWR _09506_/X sky130_fd_sc_hd__buf_1
XFILLER_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07698_ _07694_/X _07686_/X _07694_/X _13131_/X VGND VGND VPWR VPWR _07834_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09437_ _09446_/A VGND VGND VPWR VPWR _09437_/X sky130_fd_sc_hd__buf_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09368_ _09370_/A VGND VGND VPWR VPWR _09368_/X sky130_fd_sc_hd__clkbuf_1
X_08319_ _08319_/A VGND VGND VPWR VPWR _08324_/A sky130_fd_sc_hd__buf_1
X_09299_ _09309_/A VGND VGND VPWR VPWR _09312_/A sky130_fd_sc_hd__inv_2
XANTENNA_60 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_71 pc[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ _11330_/A VGND VGND VPWR VPWR _11393_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_93 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11261_ _14612_/Q _11254_/X _11130_/X _11256_/X VGND VGND VPWR VPWR _14612_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13000_ _14344_/Q VGND VGND VPWR VPWR _13000_/Y sky130_fd_sc_hd__inv_2
X_10212_ _10216_/A VGND VGND VPWR VPWR _10212_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11192_ _14630_/Q _11186_/X _11191_/X _11188_/X VGND VGND VPWR VPWR _14630_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10143_ _10143_/A VGND VGND VPWR VPWR _10164_/A sky130_fd_sc_hd__clkbuf_2
X_10074_ _10074_/A VGND VGND VPWR VPWR _10074_/X sky130_fd_sc_hd__buf_1
X_14951_ _09906_/X _14951_/D VGND VGND VPWR VPWR _14951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13902_ _15209_/Q _14537_/Q _14985_/Q _15401_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13902_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14882_ _10180_/X _14882_/D VGND VGND VPWR VPWR _14882_/Q sky130_fd_sc_hd__dfxtp_1
X_13833_ _14672_/Q _15248_/Q _14736_/Q _14704_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13833_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13764_ _15191_/Q _15159_/Q _14775_/Q _14807_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13764_/X sky130_fd_sc_hd__mux4_1
X_10976_ _10985_/A VGND VGND VPWR VPWR _10976_/X sky130_fd_sc_hd__buf_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15503_ _15591_/CLK _15503_/D VGND VGND VPWR VPWR wdata[29] sky130_fd_sc_hd__dfxtp_4
X_12715_ _12830_/A VGND VGND VPWR VPWR _12715_/X sky130_fd_sc_hd__buf_1
XFILLER_16_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13695_ _15134_/Q _15358_/Q _15326_/Q _15294_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13695_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15434_ _15601_/CLK _15434_/D VGND VGND VPWR VPWR data_address[7] sky130_fd_sc_hd__dfxtp_4
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12646_ _12634_/X _12645_/X _12450_/X _13219_/X _12383_/X VGND VGND VPWR VPWR _12646_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_62_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15365_ _08209_/X _15365_/D VGND VGND VPWR VPWR _15365_/Q sky130_fd_sc_hd__dfxtp_1
X_12577_ _12577_/A VGND VGND VPWR VPWR _12577_/X sky130_fd_sc_hd__clkbuf_4
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14316_ _15597_/CLK _14316_/D VGND VGND VPWR VPWR _14316_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11528_ _11528_/A VGND VGND VPWR VPWR _11528_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15296_ _08559_/X _15296_/D VGND VGND VPWR VPWR _15296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14247_ _14631_/Q _14599_/Q _14567_/Q _15367_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14247_/X sky130_fd_sc_hd__mux4_1
X_11459_ _11459_/A VGND VGND VPWR VPWR _11459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14178_ _14510_/Q _14478_/Q _14446_/Q _14414_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14178_/X sky130_fd_sc_hd__mux4_2
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13129_ _12590_/X _13018_/Y _13152_/S VGND VGND VPWR VPWR _13129_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08670_ _15266_/Q _08666_/X _08347_/X _08669_/X VGND VGND VPWR VPWR _15266_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07621_ _12025_/B VGND VGND VPWR VPWR _07622_/A sky130_fd_sc_hd__buf_1
XFILLER_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07552_ _15516_/Q VGND VGND VPWR VPWR _07630_/B sky130_fd_sc_hd__inv_2
XFILLER_34_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07483_ _07483_/A VGND VGND VPWR VPWR _07486_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09222_ _09227_/A VGND VGND VPWR VPWR _09222_/X sky130_fd_sc_hd__clkbuf_1
X_09153_ _09153_/A VGND VGND VPWR VPWR _09153_/X sky130_fd_sc_hd__buf_1
XFILLER_148_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08104_ _14303_/Q VGND VGND VPWR VPWR _11574_/A sky130_fd_sc_hd__inv_2
X_09084_ _09115_/A VGND VGND VPWR VPWR _09106_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08035_ _14316_/Q VGND VGND VPWR VPWR _08036_/A sky130_fd_sc_hd__buf_1
XFILLER_116_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09986_ _10354_/A VGND VGND VPWR VPWR _09986_/X sky130_fd_sc_hd__buf_1
X_08937_ _15200_/Q _08929_/X _08793_/X _08932_/X VGND VGND VPWR VPWR _15200_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08868_ _08868_/A VGND VGND VPWR VPWR _08868_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07819_ _07819_/A _07819_/B VGND VGND VPWR VPWR _07820_/C sky130_fd_sc_hd__nand2_1
XFILLER_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08799_ _09170_/A VGND VGND VPWR VPWR _08799_/X sky130_fd_sc_hd__buf_1
XFILLER_83_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10830_ _10830_/A VGND VGND VPWR VPWR _10830_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10761_ _11510_/A VGND VGND VPWR VPWR _10761_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater17 _13950_/S1 VGND VGND VPWR VPWR _13918_/S1 sky130_fd_sc_hd__clkbuf_16
Xrepeater28 _13950_/S0 VGND VGND VPWR VPWR _07542_/A sky130_fd_sc_hd__clkbuf_16
X_12500_ _12500_/A VGND VGND VPWR VPWR _12753_/A sky130_fd_sc_hd__buf_1
Xrepeater39 _07379_/A VGND VGND VPWR VPWR _14265_/S1 sky130_fd_sc_hd__clkbuf_16
XFILLER_9_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10692_ _14750_/Q _10682_/X _10691_/X _10687_/X VGND VGND VPWR VPWR _14750_/D sky130_fd_sc_hd__a22o_1
X_13480_ _13479_/X rdata[14] _13516_/S VGND VGND VPWR VPWR _13480_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12431_ _12431_/A _12431_/B VGND VGND VPWR VPWR _12432_/C sky130_fd_sc_hd__or2_1
X_15150_ _09112_/X _15150_/D VGND VGND VPWR VPWR _15150_/Q sky130_fd_sc_hd__dfxtp_1
X_12362_ _12362_/A VGND VGND VPWR VPWR _12362_/X sky130_fd_sc_hd__buf_1
XFILLER_153_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14101_ _14097_/X _14098_/X _14099_/X _14100_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14101_/X sky130_fd_sc_hd__mux4_1
X_11313_ _14596_/Q _11207_/A _11198_/X _11210_/A VGND VGND VPWR VPWR _14596_/D sky130_fd_sc_hd__a22o_1
X_12293_ _12588_/A VGND VGND VPWR VPWR _12590_/A sky130_fd_sc_hd__inv_2
X_15081_ _09389_/X _15081_/D VGND VGND VPWR VPWR _15081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11244_ _11246_/A VGND VGND VPWR VPWR _11244_/X sky130_fd_sc_hd__clkbuf_1
X_14032_ _15228_/Q _14556_/Q _15004_/Q _15420_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14032_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11175_ _11188_/A VGND VGND VPWR VPWR _11175_/X sky130_fd_sc_hd__buf_1
XFILLER_68_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10126_ _10132_/A VGND VGND VPWR VPWR _10126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14934_ _09983_/X _14934_/D VGND VGND VPWR VPWR _14934_/Q sky130_fd_sc_hd__dfxtp_1
X_10057_ _10067_/A VGND VGND VPWR VPWR _10064_/A sky130_fd_sc_hd__buf_1
XFILLER_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14865_ _10244_/X _14865_/D VGND VGND VPWR VPWR _14865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13816_ _13812_/X _13813_/X _13814_/X _13815_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13816_/X sky130_fd_sc_hd__mux4_2
XFILLER_91_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14796_ _10519_/X _14796_/D VGND VGND VPWR VPWR _14796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13747_ _14649_/Q _14617_/Q _14585_/Q _15385_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13747_/X sky130_fd_sc_hd__mux4_2
X_10959_ _10961_/A VGND VGND VPWR VPWR _10959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13678_ _14528_/Q _14496_/Q _14464_/Q _14432_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13678_/X sky130_fd_sc_hd__mux4_2
X_15417_ _07980_/X _15417_/D VGND VGND VPWR VPWR _15417_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12629_ _13319_/X _12389_/X _12475_/X _12906_/B VGND VGND VPWR VPWR _12629_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15348_ _08279_/X _15348_/D VGND VGND VPWR VPWR _15348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15279_ _08620_/X _15279_/D VGND VGND VPWR VPWR _15279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09840_ _09849_/A VGND VGND VPWR VPWR _09845_/A sky130_fd_sc_hd__buf_1
XFILLER_98_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09771_ _14991_/Q _09767_/X _09632_/X _09768_/X VGND VGND VPWR VPWR _14991_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08722_ _08722_/A VGND VGND VPWR VPWR _08722_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08653_ _15269_/Q _08647_/X _08535_/X _08648_/X VGND VGND VPWR VPWR _15269_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07604_ _07604_/A _13065_/X VGND VGND VPWR VPWR _15480_/D sky130_fd_sc_hd__and2_1
XFILLER_42_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08584_ _08644_/A VGND VGND VPWR VPWR _08605_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07535_ _15467_/Q VGND VGND VPWR VPWR _07535_/Y sky130_fd_sc_hd__inv_2
X_07466_ _07468_/A _13475_/X VGND VGND VPWR VPWR _15545_/D sky130_fd_sc_hd__and2_1
XFILLER_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09205_ _09215_/A VGND VGND VPWR VPWR _09205_/X sky130_fd_sc_hd__clkbuf_2
X_07397_ _07612_/A _13527_/X VGND VGND VPWR VPWR _15592_/D sky130_fd_sc_hd__and2_1
XFILLER_148_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09136_ _09136_/A VGND VGND VPWR VPWR _09136_/X sky130_fd_sc_hd__buf_1
XFILLER_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09067_ _15164_/Q _09065_/X _08813_/X _09066_/X VGND VGND VPWR VPWR _15164_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08018_ _15411_/Q _08014_/X _08016_/X _08017_/X VGND VGND VPWR VPWR _15411_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09969_ _10336_/A VGND VGND VPWR VPWR _09969_/X sky130_fd_sc_hd__buf_1
XFILLER_134_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12980_ _12984_/A _12980_/B _12984_/C VGND VGND VPWR VPWR _12980_/X sky130_fd_sc_hd__and3_1
XFILLER_18_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11931_ _14430_/Q _11925_/X _07958_/A _11928_/X VGND VGND VPWR VPWR _14430_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14650_ _11103_/X _14650_/D VGND VGND VPWR VPWR _14650_/Q sky130_fd_sc_hd__dfxtp_1
X_11862_ _11868_/A VGND VGND VPWR VPWR _11862_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13601_ _13600_/X _07310_/Y _13649_/S VGND VGND VPWR VPWR _13601_/X sky130_fd_sc_hd__mux2_1
X_10813_ _10813_/A VGND VGND VPWR VPWR _11553_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14581_ _11369_/X _14581_/D VGND VGND VPWR VPWR _14581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11793_ _14468_/Q _11688_/A _11567_/X _11691_/A VGND VGND VPWR VPWR _14468_/D sky130_fd_sc_hd__a22o_1
X_13532_ _13996_/X _14001_/X _13648_/S VGND VGND VPWR VPWR _13532_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10744_ _10754_/A VGND VGND VPWR VPWR _10744_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13463_ _13462_/X _13079_/X _14336_/Q VGND VGND VPWR VPWR _13463_/X sky130_fd_sc_hd__mux2_1
X_10675_ _10689_/A VGND VGND VPWR VPWR _10675_/X sky130_fd_sc_hd__clkbuf_1
X_15202_ _08922_/X _15202_/D VGND VGND VPWR VPWR _15202_/Q sky130_fd_sc_hd__dfxtp_1
X_12414_ _12414_/A VGND VGND VPWR VPWR _12414_/X sky130_fd_sc_hd__buf_1
X_13394_ _13398_/X _13395_/X _13408_/S VGND VGND VPWR VPWR _13394_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15133_ _09179_/X _15133_/D VGND VGND VPWR VPWR _15133_/Q sky130_fd_sc_hd__dfxtp_1
X_12345_ _12400_/B _13362_/X VGND VGND VPWR VPWR _12345_/X sky130_fd_sc_hd__or2_2
XFILLER_126_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15064_ _09450_/X _15064_/D VGND VGND VPWR VPWR _15064_/Q sky130_fd_sc_hd__dfxtp_1
X_12276_ _12791_/A _12199_/Y _12275_/Y _12207_/Y VGND VGND VPWR VPWR _12277_/A sky130_fd_sc_hd__a31o_1
X_14015_ _15134_/Q _15358_/Q _15326_/Q _15294_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14015_/X sky130_fd_sc_hd__mux4_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11227_ _14622_/Q _11221_/X _11087_/X _11224_/X VGND VGND VPWR VPWR _14622_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11158_ _11165_/A VGND VGND VPWR VPWR _11158_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10109_ _10111_/A VGND VGND VPWR VPWR _10109_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11089_ _11089_/A VGND VGND VPWR VPWR _11098_/A sky130_fd_sc_hd__buf_1
XFILLER_110_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14917_ _10058_/X _14917_/D VGND VGND VPWR VPWR _14917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14848_ _10307_/X _14848_/D VGND VGND VPWR VPWR _14848_/Q sky130_fd_sc_hd__dfxtp_1
X_14779_ _10579_/X _14779_/D VGND VGND VPWR VPWR _14779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07320_ _14393_/Q VGND VGND VPWR VPWR _07491_/B sky130_fd_sc_hd__inv_2
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07251_ _07252_/A _07251_/B VGND VGND VPWR VPWR _15635_/D sky130_fd_sc_hd__nor2_4
X_07182_ _07182_/A VGND VGND VPWR VPWR _07221_/A sky130_fd_sc_hd__buf_1
XFILLER_129_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09823_ _09823_/A VGND VGND VPWR VPWR _09886_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09754_ _09754_/A VGND VGND VPWR VPWR _09761_/A sky130_fd_sc_hd__buf_1
XFILLER_104_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08705_ _08705_/A VGND VGND VPWR VPWR _08710_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09685_ _09693_/A VGND VGND VPWR VPWR _09685_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08636_ _08642_/A VGND VGND VPWR VPWR _08636_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _08628_/A VGND VGND VPWR VPWR _08588_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07518_ _07569_/A VGND VGND VPWR VPWR _07568_/A sky130_fd_sc_hd__buf_1
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08498_ _10793_/A VGND VGND VPWR VPWR _09259_/A sky130_fd_sc_hd__buf_1
XFILLER_80_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07449_ _07451_/A _13439_/X VGND VGND VPWR VPWR _15557_/D sky130_fd_sc_hd__and2_1
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10460_ _10460_/A VGND VGND VPWR VPWR _10460_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09119_ _15149_/Q _09116_/X _08878_/X _09118_/X VGND VGND VPWR VPWR _15149_/D sky130_fd_sc_hd__a22o_1
X_10391_ _10398_/A VGND VGND VPWR VPWR _10391_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12130_ _12130_/A VGND VGND VPWR VPWR _12130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12061_ _12605_/A VGND VGND VPWR VPWR _12500_/A sky130_fd_sc_hd__buf_1
XFILLER_89_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11012_ _11014_/A VGND VGND VPWR VPWR _11012_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12963_ _12963_/A VGND VGND VPWR VPWR _12963_/X sky130_fd_sc_hd__buf_2
XFILLER_92_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14702_ _10909_/X _14702_/D VGND VGND VPWR VPWR _14702_/Q sky130_fd_sc_hd__dfxtp_1
X_11914_ _11926_/A VGND VGND VPWR VPWR _11915_/A sky130_fd_sc_hd__buf_1
XFILLER_73_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12894_ _12821_/X _12884_/X _12887_/X _12890_/Y _12893_/X VGND VGND VPWR VPWR _12894_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_61_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14633_ _11177_/X _14633_/D VGND VGND VPWR VPWR _14633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11845_ _11876_/A VGND VGND VPWR VPWR _11866_/A sky130_fd_sc_hd__clkbuf_2
X_14564_ _11422_/X _14564_/D VGND VGND VPWR VPWR _14564_/Q sky130_fd_sc_hd__dfxtp_1
X_11776_ _14474_/Q _11774_/X _11541_/X _11775_/X VGND VGND VPWR VPWR _14474_/D sky130_fd_sc_hd__a22o_1
XFILLER_41_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13515_ _13946_/X _13951_/X _13521_/S VGND VGND VPWR VPWR _13515_/X sky130_fd_sc_hd__mux2_1
X_10727_ _10727_/A VGND VGND VPWR VPWR _11484_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14495_ _11699_/X _14495_/D VGND VGND VPWR VPWR _14495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13446_ _13716_/X _13721_/X _14386_/Q VGND VGND VPWR VPWR _13446_/X sky130_fd_sc_hd__mux2_2
X_10658_ _10670_/A VGND VGND VPWR VPWR _10658_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13377_ _12703_/A _12662_/X _13418_/S VGND VGND VPWR VPWR _13377_/X sky130_fd_sc_hd__mux2_1
X_10589_ _10649_/A VGND VGND VPWR VPWR _10610_/A sky130_fd_sc_hd__clkbuf_2
X_15116_ _09254_/X _15116_/D VGND VGND VPWR VPWR _15116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12328_ _12727_/A VGND VGND VPWR VPWR _12328_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15047_ _09504_/X _15047_/D VGND VGND VPWR VPWR _15047_/Q sky130_fd_sc_hd__dfxtp_1
X_12259_ _12315_/A _12164_/X _12852_/A _12130_/X VGND VGND VPWR VPWR _12261_/A sky130_fd_sc_hd__o22a_1
XFILLER_123_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09470_ _09474_/A VGND VGND VPWR VPWR _09470_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08421_ _15319_/Q _08405_/X _08420_/X _08409_/X VGND VGND VPWR VPWR _15319_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08352_ _08352_/A VGND VGND VPWR VPWR _08352_/X sky130_fd_sc_hd__clkbuf_1
X_07303_ _07321_/B VGND VGND VPWR VPWR _07559_/D sky130_fd_sc_hd__buf_1
XFILLER_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08283_ _08292_/A VGND VGND VPWR VPWR _08283_/X sky130_fd_sc_hd__buf_1
XFILLER_20_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07234_ _13095_/X _07239_/B _07184_/A _07231_/A VGND VGND VPWR VPWR _15641_/D sky130_fd_sc_hd__o211a_1
X_07165_ _07271_/B _07165_/B VGND VGND VPWR VPWR _07214_/A sky130_fd_sc_hd__or2_1
XFILLER_117_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09806_ _14980_/Q _09702_/A _09691_/X _09705_/A VGND VGND VPWR VPWR _14980_/D sky130_fd_sc_hd__a22o_1
X_07998_ _08029_/A VGND VGND VPWR VPWR _07998_/X sky130_fd_sc_hd__buf_1
XFILLER_74_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09737_ _09737_/A VGND VGND VPWR VPWR _09737_/X sky130_fd_sc_hd__buf_1
XFILLER_55_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09668_ _15017_/Q _09660_/X _09667_/X _09663_/X VGND VGND VPWR VPWR _15017_/D sky130_fd_sc_hd__a22o_1
X_08619_ _15280_/Q _08617_/X _08466_/X _08618_/X VGND VGND VPWR VPWR _15280_/D sky130_fd_sc_hd__a22o_1
X_09599_ _09599_/A VGND VGND VPWR VPWR _09599_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11630_/A VGND VGND VPWR VPWR _11649_/A sky130_fd_sc_hd__clkbuf_4
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11561_ _11630_/A VGND VGND VPWR VPWR _11587_/A sky130_fd_sc_hd__buf_2
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13299_/X _13301_/X _15565_/Q VGND VGND VPWR VPWR _13300_/X sky130_fd_sc_hd__mux2_1
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10512_ _10512_/A VGND VGND VPWR VPWR _10521_/A sky130_fd_sc_hd__buf_1
X_14280_ _14948_/Q _15044_/Q _15012_/Q _15076_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14280_/X sky130_fd_sc_hd__mux4_2
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11492_ _14550_/Q _11488_/X _11489_/X _11491_/X VGND VGND VPWR VPWR _14550_/D sky130_fd_sc_hd__a22o_1
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13231_ _13232_/X _13241_/X _15562_/Q VGND VGND VPWR VPWR _13231_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10443_ _10443_/A VGND VGND VPWR VPWR _10443_/X sky130_fd_sc_hd__buf_1
X_13162_ _13161_/X _13238_/X _15565_/Q VGND VGND VPWR VPWR _13162_/X sky130_fd_sc_hd__mux2_2
XFILLER_109_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10374_ _10382_/A VGND VGND VPWR VPWR _10374_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12113_ _15580_/Q VGND VGND VPWR VPWR _12113_/X sky130_fd_sc_hd__buf_1
X_13093_ _15639_/Q data_address[4] _15667_/Q VGND VGND VPWR VPWR _13093_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12044_ _12316_/A _12337_/B VGND VGND VPWR VPWR _12333_/B sky130_fd_sc_hd__or2_1
XFILLER_2_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13995_ _15136_/Q _15360_/Q _15328_/Q _15296_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13995_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12946_ _12946_/A _12946_/B _12946_/C VGND VGND VPWR VPWR _12946_/X sky130_fd_sc_hd__or3_1
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15665_ _15666_/CLK _15665_/D VGND VGND VPWR VPWR _15665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12877_ _12228_/Y _12863_/A _12228_/A _12863_/Y VGND VGND VPWR VPWR _12877_/X sky130_fd_sc_hd__a22o_1
XANTENNA_150 rdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_161 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14616_ _11244_/X _14616_/D VGND VGND VPWR VPWR _14616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_183 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11828_ _11828_/A VGND VGND VPWR VPWR _11828_/X sky130_fd_sc_hd__clkbuf_1
X_15596_ _15601_/CLK _15596_/D VGND VGND VPWR VPWR _15596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_194 _12660_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14547_ _11500_/X _14547_/D VGND VGND VPWR VPWR _14547_/Q sky130_fd_sc_hd__dfxtp_1
X_11759_ _14479_/Q _11752_/X _11518_/X _11753_/X VGND VGND VPWR VPWR _14479_/D sky130_fd_sc_hd__a22o_1
XFILLER_146_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14478_ _11760_/X _14478_/D VGND VGND VPWR VPWR _14478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13429_ _13428_/X rdata[31] _14338_/Q VGND VGND VPWR VPWR _13429_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08970_ _08970_/A VGND VGND VPWR VPWR _08991_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07921_ _14295_/Q _14294_/Q _14298_/Q _07921_/D VGND VGND VPWR VPWR _08778_/C sky130_fd_sc_hd__or4_4
XFILLER_69_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07852_ _07852_/A VGND VGND VPWR VPWR _07852_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07783_ _07781_/X _07671_/X _07781_/X _13125_/X VGND VGND VPWR VPWR _07783_/X sky130_fd_sc_hd__o22a_1
XFILLER_56_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_48_clk _14315_/CLK VGND VGND VPWR VPWR _15648_/CLK sky130_fd_sc_hd__clkbuf_16
X_09522_ _11317_/B VGND VGND VPWR VPWR _10548_/A sky130_fd_sc_hd__buf_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09453_ _15063_/Q _09445_/X _09206_/X _09446_/X VGND VGND VPWR VPWR _15063_/D sky130_fd_sc_hd__a22o_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08404_ _08411_/A VGND VGND VPWR VPWR _08404_/X sky130_fd_sc_hd__clkbuf_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09384_ _09402_/A VGND VGND VPWR VPWR _09391_/A sky130_fd_sc_hd__buf_1
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08335_ _15332_/Q _08227_/A _08095_/X _08230_/A VGND VGND VPWR VPWR _15332_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08266_ _08270_/A VGND VGND VPWR VPWR _08266_/X sky130_fd_sc_hd__clkbuf_1
X_07217_ _07217_/A VGND VGND VPWR VPWR _07217_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08197_ _15370_/Q _08195_/X _08064_/X _08196_/X VGND VGND VPWR VPWR _15370_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07148_ _13096_/X VGND VGND VPWR VPWR _07284_/B sky130_fd_sc_hd__inv_2
XFILLER_3_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10090_ _14911_/Q _10086_/X _09944_/X _10089_/X VGND VGND VPWR VPWR _14911_/D sky130_fd_sc_hd__a22o_1
XFILLER_126_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_clk _14397_/CLK VGND VGND VPWR VPWR _15509_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12800_ _12800_/A VGND VGND VPWR VPWR _12839_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13780_ _14966_/Q _15062_/Q _15030_/Q _15094_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13780_/X sky130_fd_sc_hd__mux4_2
X_10992_ _14679_/Q _10985_/X _10728_/X _10986_/X VGND VGND VPWR VPWR _14679_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12731_ _13255_/X _12698_/X _13250_/X _12701_/X _12730_/X VGND VGND VPWR VPWR _12731_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_55_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15450_ _15662_/CLK _15450_/D VGND VGND VPWR VPWR data_address[23] sky130_fd_sc_hd__dfxtp_2
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12662_ _12662_/A VGND VGND VPWR VPWR _12662_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14401_/CLK instruction[17] VGND VGND VPWR VPWR _14401_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11613_/A VGND VGND VPWR VPWR _11613_/X sky130_fd_sc_hd__buf_1
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _08157_/X _15381_/D VGND VGND VPWR VPWR _15381_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12593_/A VGND VGND VPWR VPWR _12593_/X sky130_fd_sc_hd__buf_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _15502_/CLK _14332_/D VGND VGND VPWR VPWR _14332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ _11544_/A VGND VGND VPWR VPWR _11544_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _14661_/Q _15237_/Q _14725_/Q _14693_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14263_/X sky130_fd_sc_hd__mux4_2
X_11475_ _11475_/A VGND VGND VPWR VPWR _11475_/X sky130_fd_sc_hd__buf_1
X_13214_ _13213_/X _12851_/X _15565_/Q VGND VGND VPWR VPWR _13214_/X sky130_fd_sc_hd__mux2_1
X_10426_ _10449_/A VGND VGND VPWR VPWR _10433_/A sky130_fd_sc_hd__buf_1
XFILLER_136_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14194_ _15180_/Q _15148_/Q _14764_/Q _14796_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14194_/X sky130_fd_sc_hd__mux4_2
XFILLER_152_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13145_ _12812_/A _13002_/Y _13152_/S VGND VGND VPWR VPWR _13145_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10357_ _14838_/Q _10353_/X _10354_/X _10356_/X VGND VGND VPWR VPWR _14838_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13076_ _12674_/Y _15578_/Q _13076_/S VGND VGND VPWR VPWR _13076_/X sky130_fd_sc_hd__mux2_2
X_10288_ _10288_/A VGND VGND VPWR VPWR _10288_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12027_ _12027_/A VGND VGND VPWR VPWR _12974_/B sky130_fd_sc_hd__inv_2
XFILLER_66_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13978_ _14530_/Q _14498_/Q _14466_/Q _14434_/Q _07387_/A _14060_/S1 VGND VGND VPWR
+ VPWR _13978_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12929_ _12929_/A _12929_/B _12929_/C VGND VGND VPWR VPWR _12929_/X sky130_fd_sc_hd__or3_2
XFILLER_33_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15648_ _15648_/CLK _15648_/D VGND VGND VPWR VPWR _15648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15579_ _15579_/CLK _15579_/D VGND VGND VPWR VPWR _15579_/Q sky130_fd_sc_hd__dfxtp_1
X_08120_ _08120_/A VGND VGND VPWR VPWR _08182_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08051_ _15405_/Q _08046_/X _08048_/X _08050_/X VGND VGND VPWR VPWR _15405_/D sky130_fd_sc_hd__a22o_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08953_ _08959_/A VGND VGND VPWR VPWR _08953_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07904_ _07756_/A _15595_/Q _07756_/Y VGND VGND VPWR VPWR _07905_/A sky130_fd_sc_hd__a21oi_2
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08884_ _15212_/Q _08877_/X _08883_/X _08880_/X VGND VGND VPWR VPWR _15212_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07835_ _07835_/A VGND VGND VPWR VPWR _07835_/X sky130_fd_sc_hd__buf_1
XFILLER_110_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07766_ _13148_/X _07766_/B _07766_/C VGND VGND VPWR VPWR _07766_/X sky130_fd_sc_hd__or3_2
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09505_ _09505_/A VGND VGND VPWR VPWR _09505_/X sky130_fd_sc_hd__buf_1
XFILLER_112_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07697_ _07697_/A VGND VGND VPWR VPWR _07832_/A sky130_fd_sc_hd__inv_2
XFILLER_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09436_ _09445_/A VGND VGND VPWR VPWR _09436_/X sky130_fd_sc_hd__buf_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09367_ _15088_/Q _09365_/X _09236_/X _09366_/X VGND VGND VPWR VPWR _15088_/D sky130_fd_sc_hd__a22o_1
X_08318_ _15338_/Q _08316_/X _08064_/X _08317_/X VGND VGND VPWR VPWR _15338_/D sky130_fd_sc_hd__a22o_1
XANTENNA_50 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09298_ _09298_/A VGND VGND VPWR VPWR _09298_/X sky130_fd_sc_hd__buf_1
XANTENNA_61 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 pc[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_83 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08249_ _08251_/A VGND VGND VPWR VPWR _08249_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_94 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11260_ _11260_/A VGND VGND VPWR VPWR _11260_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10211_ _10231_/A VGND VGND VPWR VPWR _10216_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11191_ _11557_/A VGND VGND VPWR VPWR _11191_/X sky130_fd_sc_hd__buf_1
XFILLER_133_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10142_ _14894_/Q _10136_/X _10020_/X _10137_/X VGND VGND VPWR VPWR _14894_/D sky130_fd_sc_hd__a22o_1
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10073_ _10087_/A VGND VGND VPWR VPWR _10074_/A sky130_fd_sc_hd__buf_1
X_14950_ _09911_/X _14950_/D VGND VGND VPWR VPWR _14950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13901_ _13897_/X _13898_/X _13899_/X _13900_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13901_/X sky130_fd_sc_hd__mux4_1
X_14881_ _10189_/X _14881_/D VGND VGND VPWR VPWR _14881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13832_ _15216_/Q _14544_/Q _14992_/Q _15408_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13832_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13763_ _14679_/Q _15255_/Q _14743_/Q _14711_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13763_/X sky130_fd_sc_hd__mux4_2
X_10975_ _10975_/A VGND VGND VPWR VPWR _10975_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12714_ _12714_/A VGND VGND VPWR VPWR _12830_/A sky130_fd_sc_hd__buf_1
XFILLER_16_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15502_ _15502_/CLK _15502_/D VGND VGND VPWR VPWR wdata[28] sky130_fd_sc_hd__dfxtp_2
XFILLER_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13694_ _15198_/Q _15166_/Q _14782_/Q _14814_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13694_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15433_ _15648_/CLK _15433_/D VGND VGND VPWR VPWR data_address[6] sky130_fd_sc_hd__dfxtp_2
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ _12645_/A VGND VGND VPWR VPWR _12645_/X sky130_fd_sc_hd__buf_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ _08212_/X _15364_/D VGND VGND VPWR VPWR _15364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12576_ _14385_/Q _07301_/X _12565_/X _07298_/X VGND VGND VPWR VPWR _13649_/S sky130_fd_sc_hd__a31oi_4
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14315_ _14315_/CLK _14315_/D VGND VGND VPWR VPWR _14315_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _11552_/A VGND VGND VPWR VPWR _11527_/X sky130_fd_sc_hd__buf_1
X_15295_ _08562_/X _15295_/D VGND VGND VPWR VPWR _15295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14246_ _14242_/X _14243_/X _14244_/X _14245_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14246_/X sky130_fd_sc_hd__mux4_2
X_11458_ _11466_/A VGND VGND VPWR VPWR _11458_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10409_ _14826_/Q _10406_/X _10407_/X _10408_/X VGND VGND VPWR VPWR _14826_/D sky130_fd_sc_hd__a22o_1
X_14177_ _14638_/Q _14606_/Q _14574_/Q _15374_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14177_/X sky130_fd_sc_hd__mux4_2
X_11389_ _14575_/Q _11384_/X _11152_/X _11385_/X VGND VGND VPWR VPWR _14575_/D sky130_fd_sc_hd__a22o_1
XFILLER_97_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13128_ _12329_/X _13019_/Y _13152_/S VGND VGND VPWR VPWR _13128_/X sky130_fd_sc_hd__mux2_1
X_13059_ _12971_/Y _15561_/Q _13076_/S VGND VGND VPWR VPWR _13059_/X sky130_fd_sc_hd__mux2_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07620_ _15520_/Q VGND VGND VPWR VPWR _12025_/B sky130_fd_sc_hd__inv_2
XFILLER_94_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07551_ _15516_/Q _07533_/Y _15518_/Q _07534_/Y _07550_/X VGND VGND VPWR VPWR _07556_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_62_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07482_ _07482_/A _13508_/X VGND VGND VPWR VPWR _15534_/D sky130_fd_sc_hd__and2_1
XFILLER_61_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09221_ _15124_/Q _09210_/X _09220_/X _09213_/X VGND VGND VPWR VPWR _15124_/D sky130_fd_sc_hd__a22o_1
X_09152_ _09152_/A VGND VGND VPWR VPWR _09152_/X sky130_fd_sc_hd__buf_1
X_08103_ _11910_/A VGND VGND VPWR VPWR _09296_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_148_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09083_ _09083_/A VGND VGND VPWR VPWR _09083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08034_ _08034_/A VGND VGND VPWR VPWR _08034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09985_ _10011_/A VGND VGND VPWR VPWR _09985_/X sky130_fd_sc_hd__buf_1
XFILLER_115_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08936_ _08936_/A VGND VGND VPWR VPWR _08936_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08867_ _15216_/Q _08864_/X _08865_/X _08866_/X VGND VGND VPWR VPWR _15216_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07818_ _07817_/A _07816_/Y _07817_/Y _07816_/A _07810_/X VGND VGND VPWR VPWR _15452_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_45_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08798_ _08825_/A VGND VGND VPWR VPWR _08798_/X sky130_fd_sc_hd__buf_1
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07749_ _15597_/Q VGND VGND VPWR VPWR _07766_/B sky130_fd_sc_hd__inv_2
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10760_ _10760_/A VGND VGND VPWR VPWR _11510_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater18 _13740_/S1 VGND VGND VPWR VPWR _13963_/S1 sky130_fd_sc_hd__clkbuf_16
XFILLER_40_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater29 _13919_/S0 VGND VGND VPWR VPWR _13950_/S0 sky130_fd_sc_hd__buf_12
X_09419_ _15073_/Q _09410_/X _09159_/X _09413_/X VGND VGND VPWR VPWR _15073_/D sky130_fd_sc_hd__a22o_1
X_10691_ _11455_/A VGND VGND VPWR VPWR _10691_/X sky130_fd_sc_hd__buf_1
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12430_ _12357_/A _12355_/Y _12395_/Y _12394_/A _12409_/A VGND VGND VPWR VPWR _12430_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_139_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12361_ _12352_/X _12359_/X _12360_/X VGND VGND VPWR VPWR _12361_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_126_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14100_ _14966_/Q _15062_/Q _15030_/Q _15094_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14100_/X sky130_fd_sc_hd__mux4_2
XFILLER_126_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11312_ _11316_/A VGND VGND VPWR VPWR _11312_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15080_ _09391_/X _15080_/D VGND VGND VPWR VPWR _15080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12292_ _12634_/A _12117_/A _12144_/A _12289_/Y _12291_/Y VGND VGND VPWR VPWR _12292_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14031_ _14027_/X _14028_/X _14029_/X _14030_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14031_/X sky130_fd_sc_hd__mux4_1
X_11243_ _14617_/Q _11241_/X _11108_/X _11242_/X VGND VGND VPWR VPWR _14617_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11174_ _11541_/A VGND VGND VPWR VPWR _11174_/X sky130_fd_sc_hd__buf_1
XFILLER_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10125_ _10134_/A VGND VGND VPWR VPWR _10132_/A sky130_fd_sc_hd__buf_1
XFILLER_121_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14933_ _09990_/X _14933_/D VGND VGND VPWR VPWR _14933_/Q sky130_fd_sc_hd__dfxtp_1
X_10056_ _14918_/Q _10050_/X _10055_/X _10052_/X VGND VGND VPWR VPWR _14918_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14864_ _10246_/X _14864_/D VGND VGND VPWR VPWR _14864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13815_ _15122_/Q _15346_/Q _15314_/Q _15282_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13815_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14795_ _10521_/X _14795_/D VGND VGND VPWR VPWR _14795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13746_ _13742_/X _13743_/X _13744_/X _13745_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13746_/X sky130_fd_sc_hd__mux4_2
X_10958_ _14689_/Q _10951_/X _10672_/X _10954_/X VGND VGND VPWR VPWR _14689_/D sky130_fd_sc_hd__a22o_1
X_13677_ _14656_/Q _14624_/Q _14592_/Q _15392_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13677_/X sky130_fd_sc_hd__mux4_1
X_10889_ _14709_/Q _10884_/X _10740_/X _10886_/X VGND VGND VPWR VPWR _14709_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ _12946_/A _12091_/X _12611_/A _12946_/B VGND VGND VPWR VPWR _12906_/B sky130_fd_sc_hd__o22a_1
X_15416_ _07986_/X _15416_/D VGND VGND VPWR VPWR _15416_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15347_ _08281_/X _15347_/D VGND VGND VPWR VPWR _15347_/Q sky130_fd_sc_hd__dfxtp_1
X_12559_ _12561_/A _12559_/B VGND VGND VPWR VPWR _12559_/Y sky130_fd_sc_hd__nor2_1
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15278_ _08622_/X _15278_/D VGND VGND VPWR VPWR _15278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14229_ _14825_/Q _14857_/Q _14889_/Q _14921_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14229_/X sky130_fd_sc_hd__mux4_2
XFILLER_113_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09770_ _09772_/A VGND VGND VPWR VPWR _09770_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08721_ _15252_/Q _08712_/X _08442_/X _08714_/X VGND VGND VPWR VPWR _15252_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08652_ _08652_/A VGND VGND VPWR VPWR _08652_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07603_ _07604_/A _13066_/X VGND VGND VPWR VPWR _15481_/D sky130_fd_sc_hd__and2_1
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08583_ _08583_/A VGND VGND VPWR VPWR _08644_/A sky130_fd_sc_hd__buf_1
X_07534_ _13521_/S VGND VGND VPWR VPWR _07534_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07465_ _07469_/A VGND VGND VPWR VPWR _07468_/A sky130_fd_sc_hd__buf_1
XFILLER_50_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09204_ _09230_/A VGND VGND VPWR VPWR _09215_/A sky130_fd_sc_hd__buf_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07396_ _07403_/A VGND VGND VPWR VPWR _07612_/A sky130_fd_sc_hd__buf_1
X_09135_ _09135_/A VGND VGND VPWR VPWR _09135_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09066_ _09076_/A VGND VGND VPWR VPWR _09066_/X sky130_fd_sc_hd__buf_1
X_08017_ _08032_/A VGND VGND VPWR VPWR _08017_/X sky130_fd_sc_hd__buf_1
XFILLER_144_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09968_ _09976_/A VGND VGND VPWR VPWR _09968_/X sky130_fd_sc_hd__buf_1
XFILLER_58_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08919_ _09290_/A VGND VGND VPWR VPWR _08919_/X sky130_fd_sc_hd__buf_1
X_09899_ _09908_/A VGND VGND VPWR VPWR _09899_/X sky130_fd_sc_hd__buf_1
XFILLER_134_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11930_ _11932_/A VGND VGND VPWR VPWR _11930_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11861_ _11870_/A VGND VGND VPWR VPWR _11868_/A sky130_fd_sc_hd__buf_1
XFILLER_72_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13600_ _14166_/X _14171_/X _13648_/S VGND VGND VPWR VPWR _13600_/X sky130_fd_sc_hd__mux2_2
X_10812_ _10812_/A VGND VGND VPWR VPWR _10812_/X sky130_fd_sc_hd__buf_1
X_14580_ _11371_/X _14580_/D VGND VGND VPWR VPWR _14580_/Q sky130_fd_sc_hd__dfxtp_1
X_11792_ _11792_/A VGND VGND VPWR VPWR _11792_/X sky130_fd_sc_hd__clkbuf_1
X_13531_ _13530_/X _13089_/X _14337_/Q VGND VGND VPWR VPWR _13531_/X sky130_fd_sc_hd__mux2_1
X_10743_ _10773_/A VGND VGND VPWR VPWR _10754_/A sky130_fd_sc_hd__buf_1
XFILLER_41_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13462_ _13461_/X rdata[20] _13516_/S VGND VGND VPWR VPWR _13462_/X sky130_fd_sc_hd__mux2_4
X_10674_ _10674_/A VGND VGND VPWR VPWR _10689_/A sky130_fd_sc_hd__buf_2
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15201_ _08934_/X _15201_/D VGND VGND VPWR VPWR _15201_/Q sky130_fd_sc_hd__dfxtp_1
X_12413_ _12403_/X _12412_/X _12360_/X VGND VGND VPWR VPWR _12413_/Y sky130_fd_sc_hd__o21ai_2
X_13393_ _13401_/X _13394_/X _13393_/S VGND VGND VPWR VPWR _13393_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15132_ _09182_/X _15132_/D VGND VGND VPWR VPWR _15132_/Q sky130_fd_sc_hd__dfxtp_1
X_12344_ _12967_/A VGND VGND VPWR VPWR _12400_/B sky130_fd_sc_hd__buf_1
XFILLER_126_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15063_ _09452_/X _15063_/D VGND VGND VPWR VPWR _15063_/Q sky130_fd_sc_hd__dfxtp_1
X_12275_ _12275_/A _12275_/B VGND VGND VPWR VPWR _12275_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14014_ _15198_/Q _15166_/Q _14782_/Q _14814_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14014_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11226_ _11228_/A VGND VGND VPWR VPWR _11226_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11157_ _14638_/Q _11147_/X _11156_/X _11149_/X VGND VGND VPWR VPWR _14638_/D sky130_fd_sc_hd__a22o_1
XFILLER_122_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10108_ _14905_/Q _10106_/X _09973_/X _10107_/X VGND VGND VPWR VPWR _14905_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11088_ _14654_/Q _11080_/X _11087_/X _11084_/X VGND VGND VPWR VPWR _14654_/D sky130_fd_sc_hd__a22o_1
X_14916_ _10061_/X _14916_/D VGND VGND VPWR VPWR _14916_/Q sky130_fd_sc_hd__dfxtp_1
X_10039_ _10052_/A VGND VGND VPWR VPWR _10039_/X sky130_fd_sc_hd__buf_1
XFILLER_91_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14847_ _10310_/X _14847_/D VGND VGND VPWR VPWR _14847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14778_ _10581_/X _14778_/D VGND VGND VPWR VPWR _14778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13729_ _14843_/Q _14875_/Q _14907_/Q _14939_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13729_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07250_ _07252_/A _07250_/B VGND VGND VPWR VPWR _15636_/D sky130_fd_sc_hd__nor2_1
X_07181_ _13120_/X VGND VGND VPWR VPWR _07250_/B sky130_fd_sc_hd__inv_2
XFILLER_145_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09822_ _09822_/A VGND VGND VPWR VPWR _09822_/X sky130_fd_sc_hd__clkbuf_1
X_09753_ _14996_/Q _09746_/X _09607_/X _09748_/X VGND VGND VPWR VPWR _14996_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08704_ _15257_/Q _08702_/X _08408_/X _08703_/X VGND VGND VPWR VPWR _15257_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09684_ _09684_/A VGND VGND VPWR VPWR _09693_/A sky130_fd_sc_hd__buf_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08635_ _08635_/A VGND VGND VPWR VPWR _08642_/A sky130_fd_sc_hd__buf_1
XFILLER_82_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08566_ _08566_/A VGND VGND VPWR VPWR _08628_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_120_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07517_ _07517_/A _14374_/Q VGND VGND VPWR VPWR _15510_/D sky130_fd_sc_hd__and2_1
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08497_ _14312_/Q VGND VGND VPWR VPWR _10793_/A sky130_fd_sc_hd__buf_1
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07448_ _07456_/A VGND VGND VPWR VPWR _07451_/A sky130_fd_sc_hd__clkbuf_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07379_ _07379_/A VGND VGND VPWR VPWR _12569_/A sky130_fd_sc_hd__inv_2
XFILLER_136_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09118_ _09137_/A VGND VGND VPWR VPWR _09118_/X sky130_fd_sc_hd__buf_1
X_10390_ _14830_/Q _10378_/X _10389_/X _10380_/X VGND VGND VPWR VPWR _14830_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09049_ _09051_/A VGND VGND VPWR VPWR _09049_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12060_ _12448_/A VGND VGND VPWR VPWR _12605_/A sky130_fd_sc_hd__inv_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11011_ _14674_/Q _11006_/X _10756_/X _11007_/X VGND VGND VPWR VPWR _14674_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12962_ _12962_/A _12962_/B VGND VGND VPWR VPWR _12962_/Y sky130_fd_sc_hd__nor2_2
XFILLER_58_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14701_ _10912_/X _14701_/D VGND VGND VPWR VPWR _14701_/Q sky130_fd_sc_hd__dfxtp_1
X_11913_ _11923_/A VGND VGND VPWR VPWR _11926_/A sky130_fd_sc_hd__inv_2
X_12893_ _12891_/Y _12892_/Y _13354_/X _12892_/A _12681_/X VGND VGND VPWR VPWR _12893_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11844_ _11865_/A VGND VGND VPWR VPWR _11844_/X sky130_fd_sc_hd__buf_1
X_14632_ _11182_/X _14632_/D VGND VGND VPWR VPWR _14632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14563_ _11425_/X _14563_/D VGND VGND VPWR VPWR _14563_/Q sky130_fd_sc_hd__dfxtp_1
X_11775_ _11784_/A VGND VGND VPWR VPWR _11775_/X sky130_fd_sc_hd__buf_1
XFILLER_14_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10726_ _10738_/A VGND VGND VPWR VPWR _10726_/X sky130_fd_sc_hd__clkbuf_1
X_13514_ _13513_/X _13062_/X _14336_/Q VGND VGND VPWR VPWR _13514_/X sky130_fd_sc_hd__mux2_1
X_14494_ _11708_/X _14494_/D VGND VGND VPWR VPWR _14494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13445_ _13444_/X _13085_/X _14336_/Q VGND VGND VPWR VPWR _13445_/X sky130_fd_sc_hd__mux2_1
X_10657_ _10674_/A VGND VGND VPWR VPWR _10670_/A sky130_fd_sc_hd__buf_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13376_ _13378_/X _13377_/X _13415_/S VGND VGND VPWR VPWR _13376_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10588_ _10834_/A VGND VGND VPWR VPWR _10649_/A sky130_fd_sc_hd__clkbuf_2
X_12327_ _12714_/A VGND VGND VPWR VPWR _12727_/A sky130_fd_sc_hd__buf_1
X_15115_ _09258_/X _15115_/D VGND VGND VPWR VPWR _15115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15046_ _09511_/X _15046_/D VGND VGND VPWR VPWR _15046_/Q sky130_fd_sc_hd__dfxtp_1
X_12258_ _15565_/Q VGND VGND VPWR VPWR _12852_/A sky130_fd_sc_hd__inv_2
XFILLER_123_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11209_ _11222_/A VGND VGND VPWR VPWR _11210_/A sky130_fd_sc_hd__buf_1
XFILLER_141_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12189_ _12187_/X _12157_/A _12763_/A _12148_/A VGND VGND VPWR VPWR _12190_/B sky130_fd_sc_hd__o22a_1
XFILLER_68_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08420_ _09206_/A VGND VGND VPWR VPWR _08420_/X sky130_fd_sc_hd__buf_1
X_08351_ _15330_/Q _08344_/X _08347_/X _08350_/X VGND VGND VPWR VPWR _15330_/D sky130_fd_sc_hd__a22o_1
X_07302_ _14376_/Q VGND VGND VPWR VPWR _07321_/B sky130_fd_sc_hd__inv_2
XFILLER_60_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08282_ _08291_/A VGND VGND VPWR VPWR _08282_/X sky130_fd_sc_hd__buf_1
X_07233_ _07233_/A VGND VGND VPWR VPWR _07239_/B sky130_fd_sc_hd__inv_2
XFILLER_118_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07164_ _07272_/B _07217_/A VGND VGND VPWR VPWR _07165_/B sky130_fd_sc_hd__or2_2
XFILLER_117_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09805_ _09809_/A VGND VGND VPWR VPWR _09805_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07997_ _08045_/A VGND VGND VPWR VPWR _08029_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09736_ _09736_/A VGND VGND VPWR VPWR _09736_/X sky130_fd_sc_hd__buf_1
XFILLER_28_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09667_ _10411_/A VGND VGND VPWR VPWR _09667_/X sky130_fd_sc_hd__buf_1
XFILLER_131_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08618_ _08618_/A VGND VGND VPWR VPWR _08618_/X sky130_fd_sc_hd__buf_1
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09598_ _15030_/Q _09593_/X _09595_/X _09597_/X VGND VGND VPWR VPWR _15030_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08559_/A VGND VGND VPWR VPWR _08549_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ _11755_/A VGND VGND VPWR VPWR _11630_/A sky130_fd_sc_hd__buf_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10511_ _14798_/Q _10505_/X _10389_/X _10506_/X VGND VGND VPWR VPWR _14798_/D sky130_fd_sc_hd__a22o_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11491_ _11515_/A VGND VGND VPWR VPWR _11491_/X sky130_fd_sc_hd__buf_1
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13231_/X _13252_/X _15563_/Q VGND VGND VPWR VPWR _13230_/X sky130_fd_sc_hd__mux2_1
X_10442_ _10454_/A VGND VGND VPWR VPWR _10443_/A sky130_fd_sc_hd__buf_1
XFILLER_40_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13161_ _13160_/X _13200_/X _13393_/S VGND VGND VPWR VPWR _13161_/X sky130_fd_sc_hd__mux2_1
X_10373_ _10373_/A VGND VGND VPWR VPWR _10382_/A sky130_fd_sc_hd__buf_1
XFILLER_108_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12112_ _15548_/Q VGND VGND VPWR VPWR _12634_/A sky130_fd_sc_hd__inv_2
X_13092_ _15638_/Q data_address[3] _15667_/Q VGND VGND VPWR VPWR _13092_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12043_ _12979_/B VGND VGND VPWR VPWR _12337_/B sky130_fd_sc_hd__inv_2
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13994_ _15200_/Q _15168_/Q _14784_/Q _14816_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13994_/X sky130_fd_sc_hd__mux4_1
XFILLER_92_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12945_ _12643_/X _12645_/X _12908_/A _12944_/X VGND VGND VPWR VPWR _12945_/X sky130_fd_sc_hd__o22a_1
XFILLER_80_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15664_ _15666_/CLK _15664_/D VGND VGND VPWR VPWR _15664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12876_ _12670_/X _12879_/B _12384_/X VGND VGND VPWR VPWR _12876_/X sky130_fd_sc_hd__o21a_1
XANTENNA_140 rdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_151 rdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 wdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14615_ _11246_/X _14615_/D VGND VGND VPWR VPWR _14615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_184 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11827_ _14460_/Q _11825_/X _07968_/A _11826_/X VGND VGND VPWR VPWR _14460_/D sky130_fd_sc_hd__a22o_1
X_15595_ _15601_/CLK _15595_/D VGND VGND VPWR VPWR _15595_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_195 _13628_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11758_ _11762_/A VGND VGND VPWR VPWR _11758_/X sky130_fd_sc_hd__clkbuf_1
X_14546_ _11505_/X _14546_/D VGND VGND VPWR VPWR _14546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10709_ _14747_/Q _10701_/X _10708_/X _10704_/X VGND VGND VPWR VPWR _14747_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11689_ _11700_/A VGND VGND VPWR VPWR _11703_/A sky130_fd_sc_hd__inv_2
X_14477_ _11762_/X _14477_/D VGND VGND VPWR VPWR _14477_/Q sky130_fd_sc_hd__dfxtp_1
X_13428_ _13656_/X _13661_/X _13521_/S VGND VGND VPWR VPWR _13428_/X sky130_fd_sc_hd__mux2_1
X_13359_ _13358_/X _13375_/X _13393_/S VGND VGND VPWR VPWR _13359_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07920_ _07919_/Y _14296_/Q _14293_/Q _14292_/Q VGND VGND VPWR VPWR _07921_/D sky130_fd_sc_hd__o211ai_1
X_15029_ _09599_/X _15029_/D VGND VGND VPWR VPWR _15029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07851_ _07851_/A VGND VGND VPWR VPWR _07851_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07782_ _07781_/X _07674_/X _07670_/X _13127_/X VGND VGND VPWR VPWR _07804_/B sky130_fd_sc_hd__o22a_1
XFILLER_49_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09521_ _09521_/A VGND VGND VPWR VPWR _11317_/B sky130_fd_sc_hd__buf_1
XFILLER_64_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ _09454_/A VGND VGND VPWR VPWR _09452_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08403_ _15322_/Q _08387_/X _08402_/X _08391_/X VGND VGND VPWR VPWR _15322_/D sky130_fd_sc_hd__a22o_1
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09383_ _09383_/A VGND VGND VPWR VPWR _09402_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08334_ _08334_/A VGND VGND VPWR VPWR _08334_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08265_ _08285_/A VGND VGND VPWR VPWR _08270_/A sky130_fd_sc_hd__buf_2
XFILLER_137_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07216_ _07271_/B _07165_/B _07212_/X _07214_/Y VGND VGND VPWR VPWR _15651_/D sky130_fd_sc_hd__a211oi_2
X_08196_ _08205_/A VGND VGND VPWR VPWR _08196_/X sky130_fd_sc_hd__buf_1
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07147_ _13097_/X VGND VGND VPWR VPWR _07282_/B sky130_fd_sc_hd__inv_2
XFILLER_106_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09719_ _15007_/Q _09715_/X _09546_/X _09718_/X VGND VGND VPWR VPWR _15007_/D sky130_fd_sc_hd__a22o_1
X_10991_ _10993_/A VGND VGND VPWR VPWR _10991_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12730_ _12730_/A _12730_/B _12758_/C VGND VGND VPWR VPWR _12730_/X sky130_fd_sc_hd__or3_1
XFILLER_70_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12661_/A VGND VGND VPWR VPWR _12662_/A sky130_fd_sc_hd__buf_1
XFILLER_70_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11612_/A VGND VGND VPWR VPWR _11612_/X sky130_fd_sc_hd__buf_1
X_14400_ _14401_/CLK instruction[16] VGND VGND VPWR VPWR _14400_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12590_/X _12591_/X _12416_/X _13199_/X _12417_/X VGND VGND VPWR VPWR _12592_/X
+ sky130_fd_sc_hd__o32a_1
X_15380_ _08159_/X _15380_/D VGND VGND VPWR VPWR _15380_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ _15498_/CLK _14331_/D VGND VGND VPWR VPWR _14331_/Q sky130_fd_sc_hd__dfxtp_1
X_11543_ _14538_/Q _11540_/X _11541_/X _11542_/X VGND VGND VPWR VPWR _14538_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _15205_/Q _14533_/Q _14981_/Q _15397_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14262_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11474_ _11474_/A VGND VGND VPWR VPWR _11474_/X sky130_fd_sc_hd__buf_1
XFILLER_7_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13213_ _13215_/X _13257_/X _13393_/S VGND VGND VPWR VPWR _13213_/X sky130_fd_sc_hd__mux2_1
X_10425_ _10462_/A VGND VGND VPWR VPWR _10449_/A sky130_fd_sc_hd__buf_2
X_14193_ _14668_/Q _15244_/Q _14732_/Q _14700_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14193_/X sky130_fd_sc_hd__mux4_2
XFILLER_137_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13144_ _12775_/X _13003_/Y _13152_/S VGND VGND VPWR VPWR _13144_/X sky130_fd_sc_hd__mux2_2
XFILLER_3_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10356_ _10380_/A VGND VGND VPWR VPWR _10356_/X sky130_fd_sc_hd__buf_1
XFILLER_152_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13075_ _12683_/Y _15577_/Q _13076_/S VGND VGND VPWR VPWR _13075_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10287_ _14853_/Q _10280_/X _10059_/X _10281_/X VGND VGND VPWR VPWR _14853_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12026_ _12026_/A VGND VGND VPWR VPWR _12027_/A sky130_fd_sc_hd__buf_1
XFILLER_39_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13977_ _14658_/Q _14626_/Q _14594_/Q _15394_/Q _07387_/A _14060_/S1 VGND VGND VPWR
+ VPWR _13977_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12928_ _12888_/X _12926_/X _12927_/Y VGND VGND VPWR VPWR _12928_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15647_ _15647_/CLK _15647_/D VGND VGND VPWR VPWR _15647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12859_ _13305_/X VGND VGND VPWR VPWR _12859_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15578_ _15578_/CLK _15578_/D VGND VGND VPWR VPWR _15578_/Q sky130_fd_sc_hd__dfxtp_1
X_14529_ _11583_/X _14529_/D VGND VGND VPWR VPWR _14529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08050_ _08080_/A VGND VGND VPWR VPWR _08050_/X sky130_fd_sc_hd__buf_1
XFILLER_134_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08952_ _08961_/A VGND VGND VPWR VPWR _08959_/A sky130_fd_sc_hd__buf_1
X_07903_ _07900_/Y _07902_/A _07900_/A _07902_/Y _07869_/X VGND VGND VPWR VPWR _15430_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08883_ _09255_/A VGND VGND VPWR VPWR _08883_/X sky130_fd_sc_hd__buf_1
XFILLER_69_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07834_ _07834_/A VGND VGND VPWR VPWR _07834_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07765_ _07895_/A VGND VGND VPWR VPWR _07765_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09504_ _09504_/A VGND VGND VPWR VPWR _09504_/X sky130_fd_sc_hd__clkbuf_1
X_07696_ _07694_/X _13132_/X _07695_/Y VGND VGND VPWR VPWR _07697_/A sky130_fd_sc_hd__a21oi_2
XFILLER_25_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09435_ _09435_/A VGND VGND VPWR VPWR _09435_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09366_ _09366_/A VGND VGND VPWR VPWR _09366_/X sky130_fd_sc_hd__buf_1
X_08317_ _08326_/A VGND VGND VPWR VPWR _08317_/X sky130_fd_sc_hd__buf_1
XFILLER_138_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_40 data_address[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09297_ _09309_/A VGND VGND VPWR VPWR _09298_/A sky130_fd_sc_hd__buf_1
XFILLER_138_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_51 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 pc[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08248_ _15358_/Q _08241_/X _07958_/X _08244_/X VGND VGND VPWR VPWR _15358_/D sky130_fd_sc_hd__a22o_1
XANTENNA_84 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_95 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08179_ _15374_/Q _08173_/X _08042_/X _08174_/X VGND VGND VPWR VPWR _15374_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10210_ _10240_/A VGND VGND VPWR VPWR _10231_/A sky130_fd_sc_hd__buf_1
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11190_ _11190_/A VGND VGND VPWR VPWR _11190_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10141_ _10141_/A VGND VGND VPWR VPWR _10141_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10072_ _10084_/A VGND VGND VPWR VPWR _10087_/A sky130_fd_sc_hd__inv_2
XFILLER_88_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13900_ _14954_/Q _15050_/Q _15018_/Q _15082_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13900_/X sky130_fd_sc_hd__mux4_2
XFILLER_153_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14880_ _10191_/X _14880_/D VGND VGND VPWR VPWR _14880_/Q sky130_fd_sc_hd__dfxtp_1
X_13831_ _13827_/X _13828_/X _13829_/X _13830_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13831_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10974_ _14685_/Q _10964_/X _10698_/X _10967_/X VGND VGND VPWR VPWR _14685_/D sky130_fd_sc_hd__a22o_1
X_13762_ _15223_/Q _14551_/Q _14999_/Q _15415_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13762_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15501_ _15502_/CLK _15501_/D VGND VGND VPWR VPWR wdata[27] sky130_fd_sc_hd__dfxtp_2
X_12713_ _12753_/A VGND VGND VPWR VPWR _12713_/X sky130_fd_sc_hd__buf_2
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13693_ _14686_/Q _15262_/Q _14750_/Q _14718_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13693_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15432_ _15648_/CLK _15432_/D VGND VGND VPWR VPWR data_address[5] sky130_fd_sc_hd__dfxtp_1
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12644_ _12643_/X _12113_/X _12616_/X VGND VGND VPWR VPWR _12644_/Y sky130_fd_sc_hd__o21ai_2
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ _12575_/A _12575_/B VGND VGND VPWR VPWR _12575_/X sky130_fd_sc_hd__or2_1
X_15363_ _08214_/X _15363_/D VGND VGND VPWR VPWR _15363_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314_ _14381_/CLK _14314_/D VGND VGND VPWR VPWR _14314_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11526_ _11526_/A VGND VGND VPWR VPWR _11552_/A sky130_fd_sc_hd__buf_1
X_15294_ _08570_/X _15294_/D VGND VGND VPWR VPWR _15294_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11457_ _11469_/A VGND VGND VPWR VPWR _11466_/A sky130_fd_sc_hd__buf_1
X_14245_ _15111_/Q _15335_/Q _15303_/Q _15271_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14245_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10408_ _10420_/A VGND VGND VPWR VPWR _10408_/X sky130_fd_sc_hd__buf_1
X_14176_ _14172_/X _14173_/X _14174_/X _14175_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14176_/X sky130_fd_sc_hd__mux4_2
X_11388_ _11392_/A VGND VGND VPWR VPWR _11388_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13127_ _12395_/A _13020_/Y _13152_/S VGND VGND VPWR VPWR _13127_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10339_ _10339_/A VGND VGND VPWR VPWR _10339_/X sky130_fd_sc_hd__buf_1
XFILLER_152_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13058_ wdata[31] rdata[31] _13058_/S VGND VGND VPWR VPWR _14335_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12009_ _14406_/Q _12005_/X _08084_/A _12006_/X VGND VGND VPWR VPWR _14406_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_opt_3_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR clkbuf_opt_3_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07550_ _07632_/B _07541_/A _15517_/Q _07536_/Y VGND VGND VPWR VPWR _07550_/X sky130_fd_sc_hd__o22a_1
XFILLER_81_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07481_ _07482_/A _13505_/X VGND VGND VPWR VPWR _15535_/D sky130_fd_sc_hd__and2_1
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09220_ _09220_/A VGND VGND VPWR VPWR _09220_/X sky130_fd_sc_hd__buf_1
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09151_ _09167_/A VGND VGND VPWR VPWR _09152_/A sky130_fd_sc_hd__buf_1
X_08102_ _08116_/A VGND VGND VPWR VPWR _08102_/X sky130_fd_sc_hd__clkbuf_1
X_09082_ _15159_/Q _09075_/X _08834_/X _09076_/X VGND VGND VPWR VPWR _15159_/D sky130_fd_sc_hd__a22o_1
X_08033_ _15408_/Q _08029_/X _08031_/X _08032_/X VGND VGND VPWR VPWR _15408_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09984_ _10023_/A VGND VGND VPWR VPWR _10011_/A sky130_fd_sc_hd__buf_2
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08935_ _15201_/Q _08929_/X _08789_/X _08932_/X VGND VGND VPWR VPWR _15201_/D sky130_fd_sc_hd__a22o_1
XFILLER_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08866_ _08866_/A VGND VGND VPWR VPWR _08866_/X sky130_fd_sc_hd__buf_1
XFILLER_57_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07817_ _07817_/A VGND VGND VPWR VPWR _07817_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08797_ _08876_/A VGND VGND VPWR VPWR _08825_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07748_ _13148_/X VGND VGND VPWR VPWR _07748_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07679_ _07679_/A VGND VGND VPWR VPWR _07680_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater19 _07541_/A VGND VGND VPWR VPWR _13740_/S1 sky130_fd_sc_hd__clkbuf_16
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09418_ _09422_/A VGND VGND VPWR VPWR _09418_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10690_ _10690_/A VGND VGND VPWR VPWR _11455_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09349_ _09351_/A VGND VGND VPWR VPWR _09349_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12360_ _12360_/A VGND VGND VPWR VPWR _12360_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11311_ _11337_/A VGND VGND VPWR VPWR _11316_/A sky130_fd_sc_hd__buf_1
X_12291_ _12643_/A _12117_/Y _12641_/A VGND VGND VPWR VPWR _12291_/Y sky130_fd_sc_hd__o21ai_1
X_14030_ _14973_/Q _15069_/Q _15037_/Q _15101_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14030_/X sky130_fd_sc_hd__mux4_2
X_11242_ _11242_/A VGND VGND VPWR VPWR _11242_/X sky130_fd_sc_hd__buf_1
XFILLER_107_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11173_ _11186_/A VGND VGND VPWR VPWR _11173_/X sky130_fd_sc_hd__buf_1
XFILLER_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10124_ _14900_/Q _10117_/X _09995_/X _10119_/X VGND VGND VPWR VPWR _14900_/D sky130_fd_sc_hd__a22o_1
XFILLER_94_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14932_ _09994_/X _14932_/D VGND VGND VPWR VPWR _14932_/Q sky130_fd_sc_hd__dfxtp_1
X_10055_ _10423_/A VGND VGND VPWR VPWR _10055_/X sky130_fd_sc_hd__buf_1
XFILLER_0_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14863_ _10251_/X _14863_/D VGND VGND VPWR VPWR _14863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13814_ _15186_/Q _15154_/Q _14770_/Q _14802_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13814_/X sky130_fd_sc_hd__mux4_1
X_14794_ _10525_/X _14794_/D VGND VGND VPWR VPWR _14794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13745_ _15129_/Q _15353_/Q _15321_/Q _15289_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13745_/X sky130_fd_sc_hd__mux4_1
X_10957_ _10961_/A VGND VGND VPWR VPWR _10957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13676_ _13672_/X _13673_/X _13674_/X _13675_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13676_/X sky130_fd_sc_hd__mux4_2
X_10888_ _10890_/A VGND VGND VPWR VPWR _10888_/X sky130_fd_sc_hd__clkbuf_1
X_15415_ _07992_/X _15415_/D VGND VGND VPWR VPWR _15415_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ _12627_/A VGND VGND VPWR VPWR _12946_/B sky130_fd_sc_hd__buf_1
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15346_ _08286_/X _15346_/D VGND VGND VPWR VPWR _15346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12558_ data_address[1] VGND VGND VPWR VPWR _12561_/A sky130_fd_sc_hd__inv_2
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11509_ _11517_/A VGND VGND VPWR VPWR _11509_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15277_ _08625_/X _15277_/D VGND VGND VPWR VPWR _15277_/Q sky130_fd_sc_hd__dfxtp_1
X_12489_ _12860_/A _12489_/B VGND VGND VPWR VPWR _12489_/X sky130_fd_sc_hd__or2_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14228_ _14505_/Q _14473_/Q _14441_/Q _14409_/Q _14238_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14228_/X sky130_fd_sc_hd__mux4_2
XFILLER_132_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14159_ _14832_/Q _14864_/Q _14896_/Q _14928_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14159_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08720_ _08722_/A VGND VGND VPWR VPWR _08720_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08651_ _15270_/Q _08647_/X _08529_/X _08648_/X VGND VGND VPWR VPWR _15270_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07602_ _07604_/A _13067_/X VGND VGND VPWR VPWR _15482_/D sky130_fd_sc_hd__and2_1
X_08582_ _15290_/Q _08576_/X _08402_/X _08577_/X VGND VGND VPWR VPWR _15290_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07533_ _07533_/A VGND VGND VPWR VPWR _07533_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07464_ _07464_/A _13472_/X VGND VGND VPWR VPWR _15546_/D sky130_fd_sc_hd__and2_1
X_09203_ _09281_/A VGND VGND VPWR VPWR _09230_/A sky130_fd_sc_hd__clkbuf_2
X_07395_ _07420_/A VGND VGND VPWR VPWR _07403_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09134_ _15144_/Q _09126_/X _08901_/X _09127_/X VGND VGND VPWR VPWR _15144_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09065_ _09075_/A VGND VGND VPWR VPWR _09065_/X sky130_fd_sc_hd__buf_1
X_08016_ _08016_/A VGND VGND VPWR VPWR _08016_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09967_ _09993_/A VGND VGND VPWR VPWR _09976_/A sky130_fd_sc_hd__buf_1
XFILLER_131_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08918_ _08918_/A VGND VGND VPWR VPWR _08918_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09898_ _09907_/A VGND VGND VPWR VPWR _09898_/X sky130_fd_sc_hd__buf_1
X_08849_ _15220_/Q _08838_/X _08848_/X _08841_/X VGND VGND VPWR VPWR _15220_/D sky130_fd_sc_hd__a22o_1
XFILLER_45_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11860_ _14450_/Q _11856_/X _08021_/A _11857_/X VGND VGND VPWR VPWR _14450_/D sky130_fd_sc_hd__a22o_1
XFILLER_45_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10811_ _10817_/A VGND VGND VPWR VPWR _10811_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11791_ _14469_/Q _11783_/X _11564_/X _11784_/X VGND VGND VPWR VPWR _14469_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13530_ _13529_/X _14334_/D _15506_/Q VGND VGND VPWR VPWR _13530_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10742_ _10790_/A VGND VGND VPWR VPWR _10773_/A sky130_fd_sc_hd__buf_1
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10673_ _14753_/Q _10663_/X _10672_/X _10668_/X VGND VGND VPWR VPWR _14753_/D sky130_fd_sc_hd__a22o_1
X_13461_ _13766_/X _13771_/X _13521_/S VGND VGND VPWR VPWR _13461_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15200_ _08936_/X _15200_/D VGND VGND VPWR VPWR _15200_/Q sky130_fd_sc_hd__dfxtp_1
X_12412_ _12412_/A VGND VGND VPWR VPWR _12412_/X sky130_fd_sc_hd__buf_1
X_13392_ _13391_/X _13393_/X _15565_/Q VGND VGND VPWR VPWR _13392_/X sky130_fd_sc_hd__mux2_2
XFILLER_127_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15131_ _09187_/X _15131_/D VGND VGND VPWR VPWR _15131_/Q sky130_fd_sc_hd__dfxtp_1
X_12343_ _12343_/A VGND VGND VPWR VPWR _12967_/A sky130_fd_sc_hd__buf_1
X_12274_ _12274_/A VGND VGND VPWR VPWR _12754_/A sky130_fd_sc_hd__buf_1
X_15062_ _09454_/X _15062_/D VGND VGND VPWR VPWR _15062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14013_ _14686_/Q _15262_/Q _14750_/Q _14718_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14013_/X sky130_fd_sc_hd__mux4_2
X_11225_ _14623_/Q _11221_/X _11081_/X _11224_/X VGND VGND VPWR VPWR _14623_/D sky130_fd_sc_hd__a22o_1
XFILLER_122_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11156_ _11523_/A VGND VGND VPWR VPWR _11156_/X sky130_fd_sc_hd__buf_1
XFILLER_110_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10107_ _10107_/A VGND VGND VPWR VPWR _10107_/X sky130_fd_sc_hd__buf_1
XFILLER_95_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11087_ _11455_/A VGND VGND VPWR VPWR _11087_/X sky130_fd_sc_hd__buf_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14915_ _10064_/X _14915_/D VGND VGND VPWR VPWR _14915_/Q sky130_fd_sc_hd__dfxtp_1
X_10038_ _10407_/A VGND VGND VPWR VPWR _10038_/X sky130_fd_sc_hd__buf_1
XFILLER_36_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14846_ _10319_/X _14846_/D VGND VGND VPWR VPWR _14846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14777_ _10583_/X _14777_/D VGND VGND VPWR VPWR _14777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11989_ _14413_/Q _11986_/X _08048_/A _11988_/X VGND VGND VPWR VPWR _14413_/D sky130_fd_sc_hd__a22o_1
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13728_ _14523_/Q _14491_/Q _14459_/Q _14427_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13728_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13659_ _14850_/Q _14882_/Q _14914_/Q _14946_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13659_/X sky130_fd_sc_hd__mux4_1
X_07180_ _07180_/A VGND VGND VPWR VPWR _07180_/Y sky130_fd_sc_hd__inv_2
X_15329_ _08352_/X _15329_/D VGND VGND VPWR VPWR _15329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09821_ _14976_/Q _09812_/X _09539_/X _09815_/X VGND VGND VPWR VPWR _14976_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09752_ _09752_/A VGND VGND VPWR VPWR _09752_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08703_ _08703_/A VGND VGND VPWR VPWR _08703_/X sky130_fd_sc_hd__buf_1
X_09683_ _15014_/Q _09675_/X _09682_/X _09678_/X VGND VGND VPWR VPWR _15014_/D sky130_fd_sc_hd__a22o_1
X_08634_ _15275_/Q _08627_/X _08499_/X _08629_/X VGND VGND VPWR VPWR _15275_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08565_ _08587_/A VGND VGND VPWR VPWR _08565_/X sky130_fd_sc_hd__buf_1
XFILLER_81_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07516_ _07635_/A _14375_/Q VGND VGND VPWR VPWR _15511_/D sky130_fd_sc_hd__or2_1
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08496_ _08508_/A VGND VGND VPWR VPWR _08496_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07447_ _07460_/A VGND VGND VPWR VPWR _07456_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07378_ _14379_/Q VGND VGND VPWR VPWR _07510_/B sky130_fd_sc_hd__inv_2
XFILLER_129_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09117_ _09117_/A VGND VGND VPWR VPWR _09137_/A sky130_fd_sc_hd__buf_1
XFILLER_109_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09048_ _15169_/Q _09041_/X _08789_/X _09044_/X VGND VGND VPWR VPWR _15169_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11010_ _11014_/A VGND VGND VPWR VPWR _11010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12961_ _13420_/S VGND VGND VPWR VPWR _12961_/Y sky130_fd_sc_hd__inv_2
X_14700_ _10918_/X _14700_/D VGND VGND VPWR VPWR _14700_/Q sky130_fd_sc_hd__dfxtp_1
X_11912_ _11912_/A VGND VGND VPWR VPWR _11912_/X sky130_fd_sc_hd__buf_1
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12892_ _12892_/A VGND VGND VPWR VPWR _12892_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14631_ _11185_/X _14631_/D VGND VGND VPWR VPWR _14631_/Q sky130_fd_sc_hd__dfxtp_1
X_11843_ _11874_/A VGND VGND VPWR VPWR _11865_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14562_ _11427_/X _14562_/D VGND VGND VPWR VPWR _14562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11774_ _11783_/A VGND VGND VPWR VPWR _11774_/X sky130_fd_sc_hd__buf_1
XFILLER_13_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13513_ _13512_/X rdata[3] _14338_/Q VGND VGND VPWR VPWR _13513_/X sky130_fd_sc_hd__mux2_1
X_10725_ _10725_/A VGND VGND VPWR VPWR _10738_/A sky130_fd_sc_hd__clkbuf_4
X_14493_ _11710_/X _14493_/D VGND VGND VPWR VPWR _14493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13444_ _13443_/X rdata[26] _13516_/S VGND VGND VPWR VPWR _13444_/X sky130_fd_sc_hd__mux2_1
X_10656_ _14756_/Q _10550_/A _10431_/X _10553_/A VGND VGND VPWR VPWR _14756_/D sky130_fd_sc_hd__a22o_1
X_13375_ _13379_/X _13376_/X _13408_/S VGND VGND VPWR VPWR _13375_/X sky130_fd_sc_hd__mux2_1
X_10587_ _10931_/A VGND VGND VPWR VPWR _10834_/A sky130_fd_sc_hd__buf_1
XFILLER_115_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15114_ _09261_/X _15114_/D VGND VGND VPWR VPWR _15114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12326_ _12369_/A VGND VGND VPWR VPWR _12714_/A sky130_fd_sc_hd__inv_2
XFILLER_127_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15045_ _09513_/X _15045_/D VGND VGND VPWR VPWR _15045_/Q sky130_fd_sc_hd__dfxtp_1
X_12257_ _15565_/Q VGND VGND VPWR VPWR _12315_/A sky130_fd_sc_hd__buf_1
XFILLER_107_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11208_ _11219_/A VGND VGND VPWR VPWR _11222_/A sky130_fd_sc_hd__inv_2
X_12188_ _15571_/Q VGND VGND VPWR VPWR _12763_/A sky130_fd_sc_hd__inv_2
XFILLER_95_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11139_ _14642_/Q _11133_/X _11138_/X _11135_/X VGND VGND VPWR VPWR _14642_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14829_ _10391_/X _14829_/D VGND VGND VPWR VPWR _14829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08350_ _08350_/A VGND VGND VPWR VPWR _08350_/X sky130_fd_sc_hd__buf_1
X_07301_ _07301_/A VGND VGND VPWR VPWR _07301_/X sky130_fd_sc_hd__clkbuf_2
X_08281_ _08281_/A VGND VGND VPWR VPWR _08281_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07232_ _13096_/X _07231_/Y _07184_/A _07157_/B VGND VGND VPWR VPWR _15642_/D sky130_fd_sc_hd__o211a_1
XFILLER_146_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07163_ _07273_/B _07163_/B VGND VGND VPWR VPWR _07217_/A sky130_fd_sc_hd__or2_1
XFILLER_9_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09804_ _09817_/A VGND VGND VPWR VPWR _09809_/A sky130_fd_sc_hd__buf_1
XFILLER_86_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07996_ _08004_/A VGND VGND VPWR VPWR _07996_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09735_ _09741_/A VGND VGND VPWR VPWR _09735_/X sky130_fd_sc_hd__clkbuf_1
X_09666_ _10803_/A VGND VGND VPWR VPWR _10411_/A sky130_fd_sc_hd__buf_1
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08617_ _08617_/A VGND VGND VPWR VPWR _08617_/X sky130_fd_sc_hd__buf_1
XFILLER_91_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09597_ _09628_/A VGND VGND VPWR VPWR _09597_/X sky130_fd_sc_hd__buf_1
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08574_/A VGND VGND VPWR VPWR _08559_/A sky130_fd_sc_hd__buf_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ _15310_/Q _08463_/X _08478_/X _08467_/X VGND VGND VPWR VPWR _15310_/D sky130_fd_sc_hd__a22o_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10510_ _10510_/A VGND VGND VPWR VPWR _10510_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11490_ _11529_/A VGND VGND VPWR VPWR _11515_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10441_ _10451_/A VGND VGND VPWR VPWR _10454_/A sky130_fd_sc_hd__inv_2
XFILLER_148_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10372_ _14834_/Q _10366_/X _10371_/X _10368_/X VGND VGND VPWR VPWR _14834_/D sky130_fd_sc_hd__a22o_1
X_13160_ _13159_/X _13181_/X _13408_/S VGND VGND VPWR VPWR _13160_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12111_ _12089_/Y _12580_/A _12579_/A VGND VGND VPWR VPWR _12111_/Y sky130_fd_sc_hd__nand3b_2
X_13091_ _15637_/Q data_address[2] _15667_/Q VGND VGND VPWR VPWR _13091_/X sky130_fd_sc_hd__mux2_2
XFILLER_2_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12042_ _12982_/A _12037_/X _12983_/C _12040_/X _12041_/X VGND VGND VPWR VPWR _12979_/B
+ sky130_fd_sc_hd__o41a_4
XFILLER_151_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13993_ _14688_/Q _15264_/Q _14752_/Q _14720_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13993_/X sky130_fd_sc_hd__mux4_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12944_ _12652_/X _12654_/X _12909_/B _12943_/X VGND VGND VPWR VPWR _12944_/X sky130_fd_sc_hd__o22a_1
XFILLER_19_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15663_ _15663_/CLK _15663_/D VGND VGND VPWR VPWR _15663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12875_ _12875_/A _12875_/B VGND VGND VPWR VPWR _12879_/B sky130_fd_sc_hd__nor2_2
XFILLER_46_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_130 rdata[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 rdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 rdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14614_ _11252_/X _14614_/D VGND VGND VPWR VPWR _14614_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_163 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11826_ _11835_/A VGND VGND VPWR VPWR _11826_/X sky130_fd_sc_hd__buf_1
X_15594_ _15599_/CLK _15594_/D VGND VGND VPWR VPWR _15594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_174 wdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 _13630_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14545_ _11509_/X _14545_/D VGND VGND VPWR VPWR _14545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11757_ _11777_/A VGND VGND VPWR VPWR _11762_/A sky130_fd_sc_hd__clkbuf_2
X_10708_ _11467_/A VGND VGND VPWR VPWR _10708_/X sky130_fd_sc_hd__buf_1
X_14476_ _11769_/X _14476_/D VGND VGND VPWR VPWR _14476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11688_ _11688_/A VGND VGND VPWR VPWR _11688_/X sky130_fd_sc_hd__buf_1
X_13427_ _15668_/Q data_address[0] _15667_/Q VGND VGND VPWR VPWR _13427_/X sky130_fd_sc_hd__mux2_1
X_10639_ _14762_/Q _10637_/X _10407_/X _10638_/X VGND VGND VPWR VPWR _14762_/D sky130_fd_sc_hd__a22o_1
X_13358_ _13357_/X _13382_/X _13408_/S VGND VGND VPWR VPWR _13358_/X sky130_fd_sc_hd__mux2_1
X_12309_ _12316_/A _12333_/A _12337_/B _12979_/A VGND VGND VPWR VPWR _12426_/A sky130_fd_sc_hd__a211o_1
X_13289_ _13337_/X _13336_/X _13408_/S VGND VGND VPWR VPWR _13289_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15028_ _09605_/X _15028_/D VGND VGND VPWR VPWR _15028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07850_ _07848_/X _07678_/X _07849_/X VGND VGND VPWR VPWR _07851_/A sky130_fd_sc_hd__o21ai_1
XFILLER_110_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07781_ _07781_/A VGND VGND VPWR VPWR _07781_/X sky130_fd_sc_hd__buf_1
XFILLER_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09520_ _09532_/A VGND VGND VPWR VPWR _09520_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09451_ _15064_/Q _09445_/X _09200_/X _09446_/X VGND VGND VPWR VPWR _15064_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08402_ _09192_/A VGND VGND VPWR VPWR _08402_/X sky130_fd_sc_hd__buf_1
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09382_ _15083_/Q _09375_/X _09259_/X _09377_/X VGND VGND VPWR VPWR _15083_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08333_ _15333_/Q _08325_/X _08091_/X _08326_/X VGND VGND VPWR VPWR _15333_/D sky130_fd_sc_hd__a22o_1
X_08264_ _08264_/A VGND VGND VPWR VPWR _08285_/A sky130_fd_sc_hd__buf_1
XFILLER_119_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07215_ _13106_/X _07214_/Y _07209_/X _07167_/B VGND VGND VPWR VPWR _15652_/D sky130_fd_sc_hd__o211a_1
X_08195_ _08204_/A VGND VGND VPWR VPWR _08195_/X sky130_fd_sc_hd__buf_1
XFILLER_118_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07146_ _13098_/X VGND VGND VPWR VPWR _07281_/B sky130_fd_sc_hd__inv_2
XFILLER_146_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07979_ _15418_/Q _07966_/X _07978_/X _07969_/X VGND VGND VPWR VPWR _15418_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09718_ _09737_/A VGND VGND VPWR VPWR _09718_/X sky130_fd_sc_hd__buf_1
XFILLER_142_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10990_ _14680_/Q _10985_/X _10723_/X _10986_/X VGND VGND VPWR VPWR _14680_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09649_ _10399_/A VGND VGND VPWR VPWR _09649_/X sky130_fd_sc_hd__buf_1
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12660_/A VGND VGND VPWR VPWR _12660_/Y sky130_fd_sc_hd__inv_2
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11611_ _11617_/A VGND VGND VPWR VPWR _11611_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12591_/A VGND VGND VPWR VPWR _12591_/X sky130_fd_sc_hd__buf_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _15502_/CLK _14330_/D VGND VGND VPWR VPWR _14330_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _11554_/A VGND VGND VPWR VPWR _11542_/X sky130_fd_sc_hd__buf_1
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ _14257_/X _14258_/X _14259_/X _14260_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14261_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11473_ _11478_/A VGND VGND VPWR VPWR _11473_/X sky130_fd_sc_hd__clkbuf_1
X_13212_ _12610_/X _12611_/X _15561_/Q VGND VGND VPWR VPWR _13212_/X sky130_fd_sc_hd__mux2_1
X_10424_ _14822_/Q _10418_/X _10423_/X _10420_/X VGND VGND VPWR VPWR _14822_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14192_ _15212_/Q _14540_/Q _14988_/Q _15404_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14192_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13143_ _12785_/A _13004_/Y _13152_/S VGND VGND VPWR VPWR _13143_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10355_ _10395_/A VGND VGND VPWR VPWR _10380_/A sky130_fd_sc_hd__buf_2
XFILLER_98_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13074_ _12705_/Y _15576_/Q _13076_/S VGND VGND VPWR VPWR _13074_/X sky130_fd_sc_hd__mux2_1
X_10286_ _10288_/A VGND VGND VPWR VPWR _10286_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12025_ _15521_/Q _12025_/B VGND VGND VPWR VPWR _12026_/A sky130_fd_sc_hd__or2_1
XFILLER_78_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13976_ _13972_/X _13973_/X _13974_/X _13975_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _13976_/X sky130_fd_sc_hd__mux4_2
XFILLER_93_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12927_ _12927_/A VGND VGND VPWR VPWR _12927_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15646_ _15646_/CLK _15646_/D VGND VGND VPWR VPWR _15646_/Q sky130_fd_sc_hd__dfxtp_1
X_12858_ _12821_/X _12851_/X _12853_/X _12856_/Y _12857_/Y VGND VGND VPWR VPWR _12858_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11809_ _14464_/Q _11800_/X _07944_/A _11803_/X VGND VGND VPWR VPWR _14464_/D sky130_fd_sc_hd__a22o_1
X_15577_ _15578_/CLK _15577_/D VGND VGND VPWR VPWR _15577_/Q sky130_fd_sc_hd__dfxtp_1
X_12789_ _12789_/A VGND VGND VPWR VPWR _12789_/X sky130_fd_sc_hd__buf_1
XFILLER_14_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14528_ _11585_/X _14528_/D VGND VGND VPWR VPWR _14528_/Q sky130_fd_sc_hd__dfxtp_1
X_14459_ _11828_/X _14459_/D VGND VGND VPWR VPWR _14459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08951_ _15197_/Q _08943_/X _08809_/X _08946_/X VGND VGND VPWR VPWR _15197_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07902_ _07902_/A VGND VGND VPWR VPWR _07902_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08882_ _08882_/A VGND VGND VPWR VPWR _08882_/X sky130_fd_sc_hd__clkbuf_1
X_07833_ _07833_/A VGND VGND VPWR VPWR _07833_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07764_ _07754_/A _15596_/Q _07754_/Y _07900_/A VGND VGND VPWR VPWR _07895_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09503_ _15048_/Q _09496_/X _09271_/X _09497_/X VGND VGND VPWR VPWR _15048_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07695_ _07695_/A VGND VGND VPWR VPWR _07695_/Y sky130_fd_sc_hd__inv_2
X_09434_ _15069_/Q _09425_/X _09180_/X _09428_/X VGND VGND VPWR VPWR _15069_/D sky130_fd_sc_hd__a22o_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09365_ _09365_/A VGND VGND VPWR VPWR _09365_/X sky130_fd_sc_hd__buf_1
XFILLER_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08316_ _08325_/A VGND VGND VPWR VPWR _08316_/X sky130_fd_sc_hd__buf_1
XFILLER_138_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_30 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09296_ _09296_/A _09523_/B VGND VGND VPWR VPWR _09309_/A sky130_fd_sc_hd__or2_1
XANTENNA_41 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_52 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08247_ _08251_/A VGND VGND VPWR VPWR _08247_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_74 pc[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08178_ _08178_/A VGND VGND VPWR VPWR _08178_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07129_ _13115_/X VGND VGND VPWR VPWR _07256_/B sky130_fd_sc_hd__inv_2
XFILLER_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10140_ _14895_/Q _10136_/X _10016_/X _10137_/X VGND VGND VPWR VPWR _14895_/D sky130_fd_sc_hd__a22o_1
XFILLER_133_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10071_ _10071_/A VGND VGND VPWR VPWR _10071_/X sky130_fd_sc_hd__buf_1
XFILLER_153_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13830_ _14961_/Q _15057_/Q _15025_/Q _15089_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13830_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13761_ _13757_/X _13758_/X _13759_/X _13760_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13761_/X sky130_fd_sc_hd__mux4_1
X_10973_ _10975_/A VGND VGND VPWR VPWR _10973_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15500_ _15502_/CLK _15500_/D VGND VGND VPWR VPWR wdata[26] sky130_fd_sc_hd__dfxtp_1
X_12712_ _15543_/Q VGND VGND VPWR VPWR _12712_/X sky130_fd_sc_hd__clkbuf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13692_ _15230_/Q _14558_/Q _15006_/Q _15422_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13692_/X sky130_fd_sc_hd__mux4_1
X_15431_ _15669_/CLK _15431_/D VGND VGND VPWR VPWR data_address[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_43_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12643_ _12643_/A VGND VGND VPWR VPWR _12643_/X sky130_fd_sc_hd__buf_1
XFILLER_31_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15362_ _08216_/X _15362_/D VGND VGND VPWR VPWR _15362_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _12574_/A VGND VGND VPWR VPWR _12575_/A sky130_fd_sc_hd__buf_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313_ _14313_/CLK _14313_/D VGND VGND VPWR VPWR _14313_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11525_ _11532_/A VGND VGND VPWR VPWR _11525_/X sky130_fd_sc_hd__clkbuf_1
X_15293_ _08572_/X _15293_/D VGND VGND VPWR VPWR _15293_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14244_ _15175_/Q _15143_/Q _14759_/Q _14791_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14244_/X sky130_fd_sc_hd__mux4_1
X_11456_ _14558_/Q _11448_/X _11455_/X _11452_/X VGND VGND VPWR VPWR _14558_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10407_ _10407_/A VGND VGND VPWR VPWR _10407_/X sky130_fd_sc_hd__buf_1
X_14175_ _15118_/Q _15342_/Q _15310_/Q _15278_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14175_/X sky130_fd_sc_hd__mux4_1
X_11387_ _11398_/A VGND VGND VPWR VPWR _11392_/A sky130_fd_sc_hd__buf_2
XFILLER_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13126_ _12388_/X _13021_/Y _13152_/S VGND VGND VPWR VPWR _13126_/X sky130_fd_sc_hd__mux2_1
X_10338_ _10343_/A VGND VGND VPWR VPWR _10338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13057_ wdata[30] rdata[30] _13057_/S VGND VGND VPWR VPWR _14334_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10269_ _14858_/Q _10267_/X _10038_/X _10268_/X VGND VGND VPWR VPWR _14858_/D sky130_fd_sc_hd__a22o_1
XFILLER_140_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12008_ _12010_/A VGND VGND VPWR VPWR _12008_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13959_ _14820_/Q _14852_/Q _14884_/Q _14916_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13959_/X sky130_fd_sc_hd__mux4_1
X_07480_ _07482_/A _13502_/X VGND VGND VPWR VPWR _15536_/D sky130_fd_sc_hd__and2_1
XFILLER_34_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15629_ _15663_/CLK _15629_/D VGND VGND VPWR VPWR pc[24] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09150_ _09150_/A _11576_/A VGND VGND VPWR VPWR _09167_/A sky130_fd_sc_hd__or2_1
XFILLER_147_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08101_ _08118_/A VGND VGND VPWR VPWR _08116_/A sky130_fd_sc_hd__buf_1
X_09081_ _09083_/A VGND VGND VPWR VPWR _09081_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08032_ _08032_/A VGND VGND VPWR VPWR _08032_/X sky130_fd_sc_hd__buf_1
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09983_ _09990_/A VGND VGND VPWR VPWR _09983_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08934_ _08936_/A VGND VGND VPWR VPWR _08934_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08865_ _09236_/A VGND VGND VPWR VPWR _08865_/X sky130_fd_sc_hd__buf_1
XFILLER_97_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07816_ _07816_/A VGND VGND VPWR VPWR _07816_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08796_ _08796_/A VGND VGND VPWR VPWR _08876_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07747_ _07746_/A _15598_/Q _07766_/C VGND VGND VPWR VPWR _07897_/A sky130_fd_sc_hd__a21oi_2
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07678_ _13136_/X VGND VGND VPWR VPWR _07678_/X sky130_fd_sc_hd__buf_1
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09417_ _09439_/A VGND VGND VPWR VPWR _09422_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _15094_/Q _09345_/X _09211_/X _09347_/X VGND VGND VPWR VPWR _15094_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09279_ _09279_/A VGND VGND VPWR VPWR _09279_/X sky130_fd_sc_hd__buf_1
XFILLER_139_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11310_ _11310_/A VGND VGND VPWR VPWR _11337_/A sky130_fd_sc_hd__buf_2
XFILLER_126_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12290_ _12290_/A VGND VGND VPWR VPWR _12641_/A sky130_fd_sc_hd__buf_1
XFILLER_148_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11241_ _11241_/A VGND VGND VPWR VPWR _11241_/X sky130_fd_sc_hd__buf_1
XFILLER_134_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11172_ _11177_/A VGND VGND VPWR VPWR _11172_/X sky130_fd_sc_hd__clkbuf_1
X_10123_ _10123_/A VGND VGND VPWR VPWR _10123_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14931_ _09997_/X _14931_/D VGND VGND VPWR VPWR _14931_/Q sky130_fd_sc_hd__dfxtp_1
X_10054_ _10054_/A VGND VGND VPWR VPWR _10054_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14862_ _10253_/X _14862_/D VGND VGND VPWR VPWR _14862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13813_ _14674_/Q _15250_/Q _14738_/Q _14706_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13813_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14793_ _10529_/X _14793_/D VGND VGND VPWR VPWR _14793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13744_ _15193_/Q _15161_/Q _14777_/Q _14809_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13744_/X sky130_fd_sc_hd__mux4_2
X_10956_ _10956_/A VGND VGND VPWR VPWR _10961_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13675_ _15136_/Q _15360_/Q _15328_/Q _15296_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13675_/X sky130_fd_sc_hd__mux4_1
X_10887_ _14710_/Q _10884_/X _10734_/X _10886_/X VGND VGND VPWR VPWR _14710_/D sky130_fd_sc_hd__a22o_1
X_15414_ _07996_/X _15414_/D VGND VGND VPWR VPWR _15414_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ _12626_/A VGND VGND VPWR VPWR _12946_/A sky130_fd_sc_hd__buf_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15345_ _08288_/X _15345_/D VGND VGND VPWR VPWR _15345_/Q sky130_fd_sc_hd__dfxtp_1
X_12557_ _12546_/X _12556_/Y _12553_/X VGND VGND VPWR VPWR wstrobe[1] sky130_fd_sc_hd__o21a_2
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11508_ _11508_/A VGND VGND VPWR VPWR _11517_/A sky130_fd_sc_hd__buf_1
XFILLER_117_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15276_ _08631_/X _15276_/D VGND VGND VPWR VPWR _15276_/Q sky130_fd_sc_hd__dfxtp_1
X_12488_ _12770_/A _12488_/B VGND VGND VPWR VPWR _12489_/B sky130_fd_sc_hd__or2_1
XFILLER_144_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14227_ _14633_/Q _14601_/Q _14569_/Q _15369_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14227_/X sky130_fd_sc_hd__mux4_1
X_11439_ _11439_/A VGND VGND VPWR VPWR _11520_/A sky130_fd_sc_hd__buf_2
XFILLER_113_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14158_ _14512_/Q _14480_/Q _14448_/Q _14416_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14158_/X sky130_fd_sc_hd__mux4_2
XFILLER_113_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13109_ _15655_/Q data_address[20] _15667_/Q VGND VGND VPWR VPWR _13109_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14089_ _14839_/Q _14871_/Q _14903_/Q _14935_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14089_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08650_ _08652_/A VGND VGND VPWR VPWR _08650_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07601_ _07609_/A VGND VGND VPWR VPWR _07604_/A sky130_fd_sc_hd__clkbuf_1
X_08581_ _08581_/A VGND VGND VPWR VPWR _08581_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07532_ _07530_/Y _13521_/S _07531_/Y _07542_/A VGND VGND VPWR VPWR _07545_/A sky130_fd_sc_hd__o22a_1
XFILLER_34_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07463_ _07464_/A _13469_/X VGND VGND VPWR VPWR _15547_/D sky130_fd_sc_hd__and2_1
X_09202_ _09202_/A VGND VGND VPWR VPWR _09281_/A sky130_fd_sc_hd__buf_2
X_07394_ _07473_/A VGND VGND VPWR VPWR _07420_/A sky130_fd_sc_hd__buf_1
X_09133_ _09135_/A VGND VGND VPWR VPWR _09133_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09064_ _09064_/A VGND VGND VPWR VPWR _09064_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08015_ _14320_/Q VGND VGND VPWR VPWR _08016_/A sky130_fd_sc_hd__buf_1
XFILLER_78_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09966_ _10044_/A VGND VGND VPWR VPWR _09993_/A sky130_fd_sc_hd__buf_2
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08917_ _15204_/Q _08782_/A _08916_/X _08786_/A VGND VGND VPWR VPWR _15204_/D sky130_fd_sc_hd__a22o_1
X_09897_ _09897_/A VGND VGND VPWR VPWR _09897_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08848_ _09220_/A VGND VGND VPWR VPWR _08848_/X sky130_fd_sc_hd__buf_1
XFILLER_84_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08779_ _08923_/A VGND VGND VPWR VPWR _11576_/A sky130_fd_sc_hd__buf_1
XFILLER_150_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10810_ _14728_/Q _10797_/X _10809_/X _10800_/X VGND VGND VPWR VPWR _14728_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11790_ _11792_/A VGND VGND VPWR VPWR _11790_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10741_ _14741_/Q _10732_/X _10740_/X _10736_/X VGND VGND VPWR VPWR _14741_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13460_ _13459_/X _13080_/X _14336_/Q VGND VGND VPWR VPWR _13460_/X sky130_fd_sc_hd__mux2_1
X_10672_ _11437_/A VGND VGND VPWR VPWR _10672_/X sky130_fd_sc_hd__buf_1
XFILLER_9_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12411_ _12410_/A _12410_/B _12432_/B _12409_/A _12410_/Y VGND VGND VPWR VPWR _12411_/X
+ sky130_fd_sc_hd__o32a_1
X_13391_ _13390_/X _13408_/X _13393_/S VGND VGND VPWR VPWR _13391_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_20_clk _14328_/CLK VGND VGND VPWR VPWR _15592_/CLK sky130_fd_sc_hd__clkbuf_16
X_15130_ _09191_/X _15130_/D VGND VGND VPWR VPWR _15130_/Q sky130_fd_sc_hd__dfxtp_1
X_12342_ _12342_/A _12342_/B _12342_/C _12341_/X VGND VGND VPWR VPWR _12342_/X sky130_fd_sc_hd__or4b_4
XFILLER_126_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15061_ _09461_/X _15061_/D VGND VGND VPWR VPWR _15061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12273_ _12273_/A VGND VGND VPWR VPWR _12273_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14012_ _15230_/Q _14558_/Q _15006_/Q _15422_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14012_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11224_ _11242_/A VGND VGND VPWR VPWR _11224_/X sky130_fd_sc_hd__buf_1
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11155_ _11165_/A VGND VGND VPWR VPWR _11155_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10106_ _10106_/A VGND VGND VPWR VPWR _10106_/X sky130_fd_sc_hd__buf_1
X_11086_ _11086_/A VGND VGND VPWR VPWR _11086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14914_ _10068_/X _14914_/D VGND VGND VPWR VPWR _14914_/Q sky130_fd_sc_hd__dfxtp_1
X_10037_ _10050_/A VGND VGND VPWR VPWR _10037_/X sky130_fd_sc_hd__buf_1
XFILLER_91_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14845_ _10323_/X _14845_/D VGND VGND VPWR VPWR _14845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14776_ _10591_/X _14776_/D VGND VGND VPWR VPWR _14776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11988_ _12006_/A VGND VGND VPWR VPWR _11988_/X sky130_fd_sc_hd__buf_1
X_13727_ _14651_/Q _14619_/Q _14587_/Q _15387_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13727_/X sky130_fd_sc_hd__mux4_2
X_10939_ _10941_/A VGND VGND VPWR VPWR _10939_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13658_ _14530_/Q _14498_/Q _14466_/Q _14434_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13658_/X sky130_fd_sc_hd__mux4_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12609_ _12609_/A VGND VGND VPWR VPWR _12609_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13589_ _13588_/X _07310_/Y _13649_/S VGND VGND VPWR VPWR _13589_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15328_ _08358_/X _15328_/D VGND VGND VPWR VPWR _15328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15259_ _08697_/X _15259_/D VGND VGND VPWR VPWR _15259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09820_ _09822_/A VGND VGND VPWR VPWR _09820_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09751_ _14997_/Q _09746_/X _09601_/X _09748_/X VGND VGND VPWR VPWR _14997_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08702_ _08702_/A VGND VGND VPWR VPWR _08702_/X sky130_fd_sc_hd__buf_1
XFILLER_100_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09682_ _10423_/A VGND VGND VPWR VPWR _09682_/X sky130_fd_sc_hd__buf_1
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08633_ _08633_/A VGND VGND VPWR VPWR _08633_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08564_ _08626_/A VGND VGND VPWR VPWR _08587_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07515_ _07521_/A VGND VGND VPWR VPWR _07635_/A sky130_fd_sc_hd__clkbuf_1
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08495_ _08531_/A VGND VGND VPWR VPWR _08508_/A sky130_fd_sc_hd__buf_1
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07446_ _07446_/A _13436_/X VGND VGND VPWR VPWR _15558_/D sky130_fd_sc_hd__and2_1
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07377_ _07377_/A _07377_/B VGND VGND VPWR VPWR _15595_/D sky130_fd_sc_hd__nor2_1
XFILLER_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09116_ _09136_/A VGND VGND VPWR VPWR _09116_/X sky130_fd_sc_hd__buf_1
XFILLER_108_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09047_ _09051_/A VGND VGND VPWR VPWR _09047_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09949_ _09949_/A VGND VGND VPWR VPWR _09949_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12960_ _12532_/X _12952_/Y _12524_/A _12962_/B _12963_/A VGND VGND VPWR VPWR _13420_/S
+ sky130_fd_sc_hd__o221a_2
XFILLER_46_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11911_ _11923_/A VGND VGND VPWR VPWR _11912_/A sky130_fd_sc_hd__buf_1
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12891_ _13354_/X VGND VGND VPWR VPWR _12891_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14630_ _11190_/X _14630_/D VGND VGND VPWR VPWR _14630_/Q sky130_fd_sc_hd__dfxtp_1
X_11842_ _11848_/A VGND VGND VPWR VPWR _11842_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14561_ _11436_/X _14561_/D VGND VGND VPWR VPWR _14561_/Q sky130_fd_sc_hd__dfxtp_1
X_11773_ _11773_/A VGND VGND VPWR VPWR _11773_/X sky130_fd_sc_hd__clkbuf_1
X_13512_ _13936_/X _13941_/X _13521_/S VGND VGND VPWR VPWR _13512_/X sky130_fd_sc_hd__mux2_2
X_10724_ _14744_/Q _10716_/X _10723_/X _10719_/X VGND VGND VPWR VPWR _14744_/D sky130_fd_sc_hd__a22o_1
X_14492_ _11712_/X _14492_/D VGND VGND VPWR VPWR _14492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13443_ _13706_/X _13711_/X _14386_/Q VGND VGND VPWR VPWR _13443_/X sky130_fd_sc_hd__mux2_1
X_10655_ _10655_/A VGND VGND VPWR VPWR _10655_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13374_ _12138_/X _12635_/X _13418_/S VGND VGND VPWR VPWR _13374_/X sky130_fd_sc_hd__mux2_1
X_10586_ _14777_/Q _10584_/X _10340_/X _10585_/X VGND VGND VPWR VPWR _14777_/D sky130_fd_sc_hd__a22o_1
X_15113_ _09266_/X _15113_/D VGND VGND VPWR VPWR _15113_/Q sky130_fd_sc_hd__dfxtp_1
X_12325_ _12333_/B _12325_/B VGND VGND VPWR VPWR _12369_/A sky130_fd_sc_hd__or2_1
X_15044_ _09515_/X _15044_/D VGND VGND VPWR VPWR _15044_/Q sky130_fd_sc_hd__dfxtp_1
X_12256_ _15533_/Q VGND VGND VPWR VPWR _12837_/A sky130_fd_sc_hd__inv_2
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11207_ _11207_/A VGND VGND VPWR VPWR _11207_/X sky130_fd_sc_hd__buf_1
XFILLER_96_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12187_ _15571_/Q VGND VGND VPWR VPWR _12187_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11138_ _11506_/A VGND VGND VPWR VPWR _11138_/X sky130_fd_sc_hd__buf_1
XFILLER_110_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11069_ _14658_/Q _11064_/X _11065_/X _11068_/X VGND VGND VPWR VPWR _14658_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14828_ _10398_/X _14828_/D VGND VGND VPWR VPWR _14828_/Q sky130_fd_sc_hd__dfxtp_1
X_14759_ _10645_/X _14759_/D VGND VGND VPWR VPWR _14759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07300_ _14384_/Q _07505_/B VGND VGND VPWR VPWR _07301_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08280_ _15348_/Q _08272_/X _08011_/X _08274_/X VGND VGND VPWR VPWR _15348_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07231_ _07231_/A VGND VGND VPWR VPWR _07231_/Y sky130_fd_sc_hd__inv_2
X_07162_ _07276_/B _07220_/A VGND VGND VPWR VPWR _07163_/B sky130_fd_sc_hd__or2_2
XFILLER_145_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09803_ _14981_/Q _09797_/X _09687_/X _09798_/X VGND VGND VPWR VPWR _14981_/D sky130_fd_sc_hd__a22o_1
X_07995_ _15415_/Q _07981_/X _07994_/X _07984_/X VGND VGND VPWR VPWR _15415_/D sky130_fd_sc_hd__a22o_1
X_09734_ _09754_/A VGND VGND VPWR VPWR _09741_/A sky130_fd_sc_hd__buf_1
XFILLER_28_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09665_ _09665_/A VGND VGND VPWR VPWR _09665_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08616_ _08622_/A VGND VGND VPWR VPWR _08616_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09596_ _09644_/A VGND VGND VPWR VPWR _09628_/A sky130_fd_sc_hd__buf_2
XFILLER_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _08547_/A VGND VGND VPWR VPWR _08574_/A sky130_fd_sc_hd__clkbuf_4
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08478_ _09245_/A VGND VGND VPWR VPWR _08478_/X sky130_fd_sc_hd__buf_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07429_ _07429_/A VGND VGND VPWR VPWR _07432_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10440_ _10440_/A VGND VGND VPWR VPWR _10440_/X sky130_fd_sc_hd__buf_1
XFILLER_136_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10371_ _10371_/A VGND VGND VPWR VPWR _10371_/X sky130_fd_sc_hd__buf_1
XFILLER_124_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12110_ _12610_/A _12284_/B _12109_/Y VGND VGND VPWR VPWR _12579_/A sky130_fd_sc_hd__a21oi_2
X_13090_ _12537_/Y _15592_/Q _13090_/S VGND VGND VPWR VPWR _13090_/X sky130_fd_sc_hd__mux2_2
XFILLER_124_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12041_ _07637_/B _12040_/X _07123_/A VGND VGND VPWR VPWR _12041_/X sky130_fd_sc_hd__o21a_1
XFILLER_105_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13992_ _15232_/Q _14560_/Q _15008_/Q _15424_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13992_/X sky130_fd_sc_hd__mux4_1
X_12943_ _12132_/X _12676_/A _12908_/B _12666_/X _12668_/X VGND VGND VPWR VPWR _12943_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_34_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15662_ _15662_/CLK _15662_/D VGND VGND VPWR VPWR _15662_/Q sky130_fd_sc_hd__dfxtp_1
X_12874_ _12874_/A _12929_/B VGND VGND VPWR VPWR _12874_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_120 rdata[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_131 rdata[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_142 rdata[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_153 rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14613_ _11258_/X _14613_/D VGND VGND VPWR VPWR _14613_/Q sky130_fd_sc_hd__dfxtp_1
X_11825_ _11834_/A VGND VGND VPWR VPWR _11825_/X sky130_fd_sc_hd__buf_1
X_15593_ _15599_/CLK _15593_/D VGND VGND VPWR VPWR _15593_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_164 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_175 wdata[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_186 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14544_ _11512_/X _14544_/D VGND VGND VPWR VPWR _14544_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_197 _13626_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11756_ _11820_/A VGND VGND VPWR VPWR _11777_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10707_ _10707_/A VGND VGND VPWR VPWR _11467_/A sky130_fd_sc_hd__buf_1
X_14475_ _11771_/X _14475_/D VGND VGND VPWR VPWR _14475_/Q sky130_fd_sc_hd__dfxtp_1
X_11687_ _11700_/A VGND VGND VPWR VPWR _11688_/A sky130_fd_sc_hd__buf_1
X_13426_ _15669_/Q data_address[1] _15667_/Q VGND VGND VPWR VPWR _13426_/X sky130_fd_sc_hd__mux2_1
X_10638_ _10647_/A VGND VGND VPWR VPWR _10638_/X sky130_fd_sc_hd__buf_1
XFILLER_127_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13357_ _13356_/X _13385_/X _13415_/S VGND VGND VPWR VPWR _13357_/X sky130_fd_sc_hd__mux2_1
X_10569_ _10578_/A VGND VGND VPWR VPWR _10574_/A sky130_fd_sc_hd__buf_1
XFILLER_115_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12308_ _12337_/A _12338_/A VGND VGND VPWR VPWR _12979_/A sky130_fd_sc_hd__and2_2
X_13288_ _12812_/A _12820_/X _15561_/Q VGND VGND VPWR VPWR _13288_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15027_ _09609_/X _15027_/D VGND VGND VPWR VPWR _15027_/Q sky130_fd_sc_hd__dfxtp_1
X_12239_ _15536_/Q _12239_/B VGND VGND VPWR VPWR _12239_/X sky130_fd_sc_hd__or2_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07780_ _07819_/B _07817_/A _07819_/A VGND VGND VPWR VPWR _07804_/A sky130_fd_sc_hd__or3_1
XFILLER_96_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09450_ _09454_/A VGND VGND VPWR VPWR _09450_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08401_ _10712_/A VGND VGND VPWR VPWR _09192_/A sky130_fd_sc_hd__buf_1
X_09381_ _09381_/A VGND VGND VPWR VPWR _09381_/X sky130_fd_sc_hd__clkbuf_1
X_08332_ _08334_/A VGND VGND VPWR VPWR _08332_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08263_ _15353_/Q _08261_/X _07983_/X _08262_/X VGND VGND VPWR VPWR _15353_/D sky130_fd_sc_hd__a22o_1
X_07214_ _07214_/A VGND VGND VPWR VPWR _07214_/Y sky130_fd_sc_hd__inv_2
X_08194_ _08200_/A VGND VGND VPWR VPWR _08194_/X sky130_fd_sc_hd__clkbuf_1
X_07145_ _13099_/X VGND VGND VPWR VPWR _07280_/B sky130_fd_sc_hd__inv_2
XFILLER_106_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07978_ _07978_/A VGND VGND VPWR VPWR _07978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09717_ _09778_/A VGND VGND VPWR VPWR _09737_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09648_ _10787_/A VGND VGND VPWR VPWR _10399_/A sky130_fd_sc_hd__buf_1
XFILLER_83_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _10340_/A VGND VGND VPWR VPWR _09579_/X sky130_fd_sc_hd__buf_1
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11610_ _11619_/A VGND VGND VPWR VPWR _11617_/A sky130_fd_sc_hd__buf_1
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12590_ _12590_/A VGND VGND VPWR VPWR _12590_/X sky130_fd_sc_hd__buf_4
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _11541_/A VGND VGND VPWR VPWR _11541_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ _14950_/Q _15046_/Q _15014_/Q _15078_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14260_/X sky130_fd_sc_hd__mux4_2
XFILLER_11_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ _14554_/Q _11462_/X _11471_/X _11464_/X VGND VGND VPWR VPWR _14554_/D sky130_fd_sc_hd__a22o_1
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13211_ _13212_/X _13222_/X _15562_/Q VGND VGND VPWR VPWR _13211_/X sky130_fd_sc_hd__mux2_1
X_10423_ _10423_/A VGND VGND VPWR VPWR _10423_/X sky130_fd_sc_hd__buf_1
X_14191_ _14187_/X _14188_/X _14189_/X _14190_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14191_/X sky130_fd_sc_hd__mux4_2
XFILLER_109_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13142_ _12762_/X _13005_/Y _13152_/S VGND VGND VPWR VPWR _13142_/X sky130_fd_sc_hd__mux2_1
X_10354_ _10354_/A VGND VGND VPWR VPWR _10354_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13073_ _12719_/Y _15575_/Q _13076_/S VGND VGND VPWR VPWR _13073_/X sky130_fd_sc_hd__mux2_1
X_10285_ _14854_/Q _10280_/X _10055_/X _10281_/X VGND VGND VPWR VPWR _14854_/D sky130_fd_sc_hd__a22o_1
XFILLER_151_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12024_ _12024_/A VGND VGND VPWR VPWR _12024_/X sky130_fd_sc_hd__buf_1
XFILLER_104_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13975_ _15138_/Q _15362_/Q _15330_/Q _15298_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13975_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12926_ _12926_/A _12926_/B VGND VGND VPWR VPWR _12926_/X sky130_fd_sc_hd__or2_1
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15645_ _15647_/CLK _15645_/D VGND VGND VPWR VPWR _15645_/Q sky130_fd_sc_hd__dfxtp_1
X_12857_ _12839_/A _12839_/B _12428_/A _12839_/Y VGND VGND VPWR VPWR _12857_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11808_ _11818_/A VGND VGND VPWR VPWR _11808_/X sky130_fd_sc_hd__clkbuf_1
X_15576_ _15576_/CLK _15576_/D VGND VGND VPWR VPWR _15576_/Q sky130_fd_sc_hd__dfxtp_1
X_12788_ _12788_/A VGND VGND VPWR VPWR _12788_/X sky130_fd_sc_hd__buf_1
XFILLER_14_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11739_ _14485_/Q _11733_/X _11494_/X _11735_/X VGND VGND VPWR VPWR _14485_/D sky130_fd_sc_hd__a22o_1
X_14527_ _11588_/X _14527_/D VGND VGND VPWR VPWR _14527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14458_ _11831_/X _14458_/D VGND VGND VPWR VPWR _14458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13409_ _13411_/X _13410_/X _13415_/S VGND VGND VPWR VPWR _13409_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14389_ _14393_/CLK instruction[26] VGND VGND VPWR VPWR _14389_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08950_ _08950_/A VGND VGND VPWR VPWR _08950_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07901_ _07754_/A _15596_/Q _07754_/Y VGND VGND VPWR VPWR _07902_/A sky130_fd_sc_hd__a21oi_2
XFILLER_69_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08881_ _15213_/Q _08877_/X _08878_/X _08880_/X VGND VGND VPWR VPWR _15213_/D sky130_fd_sc_hd__a22o_1
XFILLER_111_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07832_ _07832_/A _07832_/B VGND VGND VPWR VPWR _07833_/A sky130_fd_sc_hd__or2_1
XFILLER_57_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07763_ _07756_/A _15595_/Q _07756_/Y _07762_/Y VGND VGND VPWR VPWR _07900_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09502_ _09504_/A VGND VGND VPWR VPWR _09502_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07694_ _07701_/A VGND VGND VPWR VPWR _07694_/X sky130_fd_sc_hd__buf_1
XFILLER_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09433_ _09435_/A VGND VGND VPWR VPWR _09433_/X sky130_fd_sc_hd__clkbuf_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ _09370_/A VGND VGND VPWR VPWR _09364_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08315_ _08315_/A VGND VGND VPWR VPWR _08315_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 data_address[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09295_ _09810_/B VGND VGND VPWR VPWR _09523_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA_31 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_42 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 instruction[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08246_ _08255_/A VGND VGND VPWR VPWR _08251_/A sky130_fd_sc_hd__buf_1
XANTENNA_64 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_86 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08177_ _15375_/Q _08173_/X _08036_/X _08174_/X VGND VGND VPWR VPWR _15375_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07128_ _13116_/X VGND VGND VPWR VPWR _07255_/B sky130_fd_sc_hd__inv_2
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10070_ _10084_/A VGND VGND VPWR VPWR _10071_/A sky130_fd_sc_hd__buf_1
XFILLER_102_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13760_ _14968_/Q _15064_/Q _15032_/Q _15096_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13760_/X sky130_fd_sc_hd__mux4_1
X_10972_ _14686_/Q _10964_/X _10691_/X _10967_/X VGND VGND VPWR VPWR _14686_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12711_ _12708_/X _12709_/X _12677_/X _13249_/X _12710_/X VGND VGND VPWR VPWR _12711_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13691_ _13687_/X _13688_/X _13689_/X _13690_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13691_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15430_ _15668_/CLK _15430_/D VGND VGND VPWR VPWR data_address[3] sky130_fd_sc_hd__dfxtp_4
X_12642_ _12641_/A _12641_/B _12640_/Y _12640_/A _12641_/Y VGND VGND VPWR VPWR _12642_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ _08234_/X _15361_/D VGND VGND VPWR VPWR _15361_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ _12573_/A _12575_/B VGND VGND VPWR VPWR _12573_/X sky130_fd_sc_hd__or2_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11524_ _14542_/Q _11513_/X _11523_/X _11515_/X VGND VGND VPWR VPWR _14542_/D sky130_fd_sc_hd__a22o_1
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14312_ _14381_/CLK _14312_/D VGND VGND VPWR VPWR _14312_/Q sky130_fd_sc_hd__dfxtp_1
X_15292_ _08575_/X _15292_/D VGND VGND VPWR VPWR _15292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _14663_/Q _15239_/Q _14727_/Q _14695_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14243_/X sky130_fd_sc_hd__mux4_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11455_ _11455_/A VGND VGND VPWR VPWR _11455_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10406_ _10418_/A VGND VGND VPWR VPWR _10406_/X sky130_fd_sc_hd__buf_1
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14174_ _15182_/Q _15150_/Q _14766_/Q _14798_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14174_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11386_ _14576_/Q _11384_/X _11148_/X _11385_/X VGND VGND VPWR VPWR _14576_/D sky130_fd_sc_hd__a22o_1
XFILLER_98_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13125_ _12415_/X _13022_/Y _13152_/S VGND VGND VPWR VPWR _13125_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10337_ _14842_/Q _10327_/X _10336_/X _10329_/X VGND VGND VPWR VPWR _14842_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13056_ wdata[29] rdata[29] _13057_/S VGND VGND VPWR VPWR _14333_/D sky130_fd_sc_hd__mux2_1
X_10268_ _10281_/A VGND VGND VPWR VPWR _10268_/X sky130_fd_sc_hd__buf_1
X_12007_ _14407_/Q _12005_/X _08079_/A _12006_/X VGND VGND VPWR VPWR _14407_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10199_ _10218_/A VGND VGND VPWR VPWR _10199_/X sky130_fd_sc_hd__buf_1
XFILLER_78_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13958_ _14500_/Q _14468_/Q _14436_/Q _14404_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13958_/X sky130_fd_sc_hd__mux4_2
XFILLER_34_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12909_ _12909_/A _12909_/B _12909_/C _12909_/D VGND VGND VPWR VPWR _12959_/D sky130_fd_sc_hd__or4_4
XFILLER_62_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13889_ _14827_/Q _14859_/Q _14891_/Q _14923_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13889_/X sky130_fd_sc_hd__mux4_1
X_15628_ _15666_/CLK _15628_/D VGND VGND VPWR VPWR pc[23] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15559_ _15590_/CLK _15559_/D VGND VGND VPWR VPWR _15559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08100_ _15395_/Q _07927_/A _08099_/X _07932_/A VGND VGND VPWR VPWR _15395_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09080_ _15160_/Q _09075_/X _08830_/X _09076_/X VGND VGND VPWR VPWR _15160_/D sky130_fd_sc_hd__a22o_1
X_08031_ _08031_/A VGND VGND VPWR VPWR _08031_/X sky130_fd_sc_hd__clkbuf_2
X_09982_ _14935_/Q _09972_/X _09981_/X _09974_/X VGND VGND VPWR VPWR _14935_/D sky130_fd_sc_hd__a22o_1
XFILLER_107_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08933_ _15202_/Q _08929_/X _08783_/X _08932_/X VGND VGND VPWR VPWR _15202_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08864_ _08864_/A VGND VGND VPWR VPWR _08864_/X sky130_fd_sc_hd__buf_1
XFILLER_97_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07815_ _07813_/X _07674_/X _07820_/B VGND VGND VPWR VPWR _07816_/A sky130_fd_sc_hd__o21ai_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08795_ _08804_/A VGND VGND VPWR VPWR _08795_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07746_ _07746_/A _15598_/Q VGND VGND VPWR VPWR _07766_/C sky130_fd_sc_hd__nor2_1
XFILLER_44_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07677_ _07675_/X _13127_/X _07675_/X _13127_/X VGND VGND VPWR VPWR _07817_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09416_ _09478_/A VGND VGND VPWR VPWR _09439_/A sky130_fd_sc_hd__buf_2
XFILLER_25_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09347_ _09366_/A VGND VGND VPWR VPWR _09347_/X sky130_fd_sc_hd__buf_1
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09278_ _09278_/A VGND VGND VPWR VPWR _09278_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08229_ _08242_/A VGND VGND VPWR VPWR _08230_/A sky130_fd_sc_hd__buf_1
XFILLER_138_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11240_ _11246_/A VGND VGND VPWR VPWR _11240_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11171_ _14635_/Q _11160_/X _11170_/X _11163_/X VGND VGND VPWR VPWR _14635_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10122_ _14901_/Q _10117_/X _09991_/X _10119_/X VGND VGND VPWR VPWR _14901_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14930_ _10002_/X _14930_/D VGND VGND VPWR VPWR _14930_/Q sky130_fd_sc_hd__dfxtp_1
X_10053_ _14919_/Q _10050_/X _10051_/X _10052_/X VGND VGND VPWR VPWR _14919_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14861_ _10255_/X _14861_/D VGND VGND VPWR VPWR _14861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13812_ _15218_/Q _14546_/Q _14994_/Q _15410_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13812_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14792_ _10531_/X _14792_/D VGND VGND VPWR VPWR _14792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13743_ _14681_/Q _15257_/Q _14745_/Q _14713_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13743_/X sky130_fd_sc_hd__mux4_2
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10955_ _14690_/Q _10951_/X _10665_/X _10954_/X VGND VGND VPWR VPWR _14690_/D sky130_fd_sc_hd__a22o_1
XFILLER_44_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10886_ _10905_/A VGND VGND VPWR VPWR _10886_/X sky130_fd_sc_hd__buf_1
X_13674_ _15200_/Q _15168_/Q _14784_/Q _14816_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13674_/X sky130_fd_sc_hd__mux4_1
X_15413_ _08004_/X _15413_/D VGND VGND VPWR VPWR _15413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12625_ _12625_/A _12625_/B VGND VGND VPWR VPWR _12625_/X sky130_fd_sc_hd__or2_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12556_ _12556_/A _12561_/B VGND VGND VPWR VPWR _12556_/Y sky130_fd_sc_hd__nor2_1
X_15344_ _08290_/X _15344_/D VGND VGND VPWR VPWR _15344_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11507_ _14546_/Q _11501_/X _11506_/X _11503_/X VGND VGND VPWR VPWR _14546_/D sky130_fd_sc_hd__a22o_1
XFILLER_145_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ _12796_/A _13396_/X VGND VGND VPWR VPWR _12488_/B sky130_fd_sc_hd__or2_1
X_15275_ _08633_/X _15275_/D VGND VGND VPWR VPWR _15275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11438_ _14561_/Q _11430_/X _11437_/X _11434_/X VGND VGND VPWR VPWR _14561_/D sky130_fd_sc_hd__a22o_1
X_14226_ _14222_/X _14223_/X _14224_/X _14225_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14226_/X sky130_fd_sc_hd__mux4_2
XFILLER_153_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14157_ _14640_/Q _14608_/Q _14576_/Q _15376_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14157_/X sky130_fd_sc_hd__mux4_2
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11369_ _11373_/A VGND VGND VPWR VPWR _11369_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13108_ _15654_/Q data_address[19] _15667_/Q VGND VGND VPWR VPWR _13108_/X sky130_fd_sc_hd__mux2_1
X_14088_ _14519_/Q _14487_/Q _14455_/Q _14423_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14088_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13039_ wdata[12] rdata[12] ren VGND VGND VPWR VPWR _14316_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07600_ _07809_/A VGND VGND VPWR VPWR _07609_/A sky130_fd_sc_hd__buf_1
XFILLER_54_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08580_ _15291_/Q _08576_/X _08396_/X _08577_/X VGND VGND VPWR VPWR _15291_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07531_ _15466_/Q VGND VGND VPWR VPWR _07531_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07462_ _07464_/A _13466_/X VGND VGND VPWR VPWR _15548_/D sky130_fd_sc_hd__and2_1
XFILLER_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09201_ _15128_/Q _09195_/X _09200_/X _09197_/X VGND VGND VPWR VPWR _15128_/D sky130_fd_sc_hd__a22o_1
X_07393_ _07586_/A VGND VGND VPWR VPWR _07473_/A sky130_fd_sc_hd__buf_1
X_09132_ _15145_/Q _09126_/X _08895_/X _09127_/X VGND VGND VPWR VPWR _15145_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09063_ _15165_/Q _09054_/X _08809_/X _09057_/X VGND VGND VPWR VPWR _15165_/D sky130_fd_sc_hd__a22o_1
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08014_ _08029_/A VGND VGND VPWR VPWR _08014_/X sky130_fd_sc_hd__buf_1
XFILLER_151_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09965_ _10173_/A VGND VGND VPWR VPWR _10044_/A sky130_fd_sc_hd__clkbuf_2
X_08916_ _09287_/A VGND VGND VPWR VPWR _08916_/X sky130_fd_sc_hd__buf_1
XFILLER_134_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09896_ _14955_/Q _09887_/X _09657_/X _09889_/X VGND VGND VPWR VPWR _14955_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08847_ _08855_/A VGND VGND VPWR VPWR _08847_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08778_ _14299_/Q _14300_/Q _08778_/C VGND VGND VPWR VPWR _08923_/A sky130_fd_sc_hd__or3_1
X_07729_ _15601_/Q VGND VGND VPWR VPWR _07730_/B sky130_fd_sc_hd__inv_2
XFILLER_150_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10740_ _11494_/A VGND VGND VPWR VPWR _10740_/X sky130_fd_sc_hd__buf_1
X_10671_ _10671_/A VGND VGND VPWR VPWR _11437_/A sky130_fd_sc_hd__buf_1
XFILLER_9_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12410_ _12410_/A _12410_/B VGND VGND VPWR VPWR _12410_/Y sky130_fd_sc_hd__nor2_1
X_13390_ _13389_/X _13415_/X _13408_/S VGND VGND VPWR VPWR _13390_/X sky130_fd_sc_hd__mux2_1
X_12341_ _12329_/X _12330_/X _12336_/X _13195_/X _12493_/A VGND VGND VPWR VPWR _12341_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_138_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15060_ _09463_/X _15060_/D VGND VGND VPWR VPWR _15060_/Q sky130_fd_sc_hd__dfxtp_1
X_12272_ _15541_/Q _12168_/Y _12271_/Y _12175_/Y VGND VGND VPWR VPWR _12273_/A sky130_fd_sc_hd__a31o_1
XFILLER_107_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14011_ _14007_/X _14008_/X _14009_/X _14010_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14011_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11223_ _11285_/A VGND VGND VPWR VPWR _11242_/A sky130_fd_sc_hd__buf_2
XFILLER_122_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11154_ _11168_/A VGND VGND VPWR VPWR _11165_/A sky130_fd_sc_hd__buf_2
XFILLER_150_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10105_ _10111_/A VGND VGND VPWR VPWR _10105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11085_ _14655_/Q _11080_/X _11081_/X _11084_/X VGND VGND VPWR VPWR _14655_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14913_ _10076_/X _14913_/D VGND VGND VPWR VPWR _14913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10036_ _10041_/A VGND VGND VPWR VPWR _10036_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14844_ _10326_/X _14844_/D VGND VGND VPWR VPWR _14844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14775_ _10593_/X _14775_/D VGND VGND VPWR VPWR _14775_/Q sky130_fd_sc_hd__dfxtp_1
X_11987_ _11987_/A VGND VGND VPWR VPWR _12006_/A sky130_fd_sc_hd__clkbuf_2
X_13726_ _13722_/X _13723_/X _13724_/X _13725_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13726_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10938_ _14695_/Q _10936_/X _10814_/X _10937_/X VGND VGND VPWR VPWR _14695_/D sky130_fd_sc_hd__a22o_1
X_10869_ _10869_/A VGND VGND VPWR VPWR _10869_/X sky130_fd_sc_hd__clkbuf_1
X_13657_ _14658_/Q _14626_/Q _14594_/Q _15394_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13657_/X sky130_fd_sc_hd__mux4_2
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12608_ _12535_/X _12586_/B _12598_/Y _12601_/X _12607_/X VGND VGND VPWR VPWR _12609_/A
+ sky130_fd_sc_hd__o311a_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13588_ _14136_/X _14141_/X _13648_/S VGND VGND VPWR VPWR _13588_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15327_ _08363_/X _15327_/D VGND VGND VPWR VPWR _15327_/Q sky130_fd_sc_hd__dfxtp_1
X_12539_ _12538_/X _15459_/Q _15460_/Q VGND VGND VPWR VPWR _12541_/B sky130_fd_sc_hd__and3b_1
XFILLER_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15258_ _08699_/X _15258_/D VGND VGND VPWR VPWR _15258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14209_ _14827_/Q _14859_/Q _14891_/Q _14923_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14209_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15189_ _08978_/X _15189_/D VGND VGND VPWR VPWR _15189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09750_ _09752_/A VGND VGND VPWR VPWR _09750_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08701_ _08701_/A VGND VGND VPWR VPWR _08701_/X sky130_fd_sc_hd__clkbuf_1
X_09681_ _10818_/A VGND VGND VPWR VPWR _10423_/A sky130_fd_sc_hd__buf_1
XFILLER_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08632_ _15276_/Q _08627_/X _08492_/X _08629_/X VGND VGND VPWR VPWR _15276_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08563_ _08563_/A VGND VGND VPWR VPWR _08626_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07514_ _07514_/A _07559_/D VGND VGND VPWR VPWR _15512_/D sky130_fd_sc_hd__nor2_1
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08494_ _08547_/A VGND VGND VPWR VPWR _08531_/A sky130_fd_sc_hd__buf_1
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07445_ _07446_/A _13433_/X VGND VGND VPWR VPWR _15559_/D sky130_fd_sc_hd__and2_1
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07376_ _07377_/B VGND VGND VPWR VPWR _07376_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09115_ _09115_/A VGND VGND VPWR VPWR _09136_/A sky130_fd_sc_hd__buf_1
X_09046_ _09059_/A VGND VGND VPWR VPWR _09051_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_117_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09948_ _14943_/Q _09943_/X _09944_/X _09947_/X VGND VGND VPWR VPWR _14943_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09879_ _14960_/Q _09877_/X _09627_/X _09878_/X VGND VGND VPWR VPWR _14960_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11910_ _11910_/A _11910_/B VGND VGND VPWR VPWR _11923_/A sky130_fd_sc_hd__or2_2
X_12890_ _12796_/A _12888_/X _12829_/X _12889_/X VGND VGND VPWR VPWR _12890_/Y sky130_fd_sc_hd__o22ai_4
X_11841_ _14455_/Q _11834_/X _07994_/A _11835_/X VGND VGND VPWR VPWR _14455_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11772_ _14475_/Q _11764_/X _11537_/X _11766_/X VGND VGND VPWR VPWR _14475_/D sky130_fd_sc_hd__a22o_1
X_14560_ _11442_/X _14560_/D VGND VGND VPWR VPWR _14560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10723_ _11479_/A VGND VGND VPWR VPWR _10723_/X sky130_fd_sc_hd__buf_1
X_13511_ _13510_/X _13063_/X _14336_/Q VGND VGND VPWR VPWR _13511_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14491_ _11717_/X _14491_/D VGND VGND VPWR VPWR _14491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13442_ _13441_/X _13086_/X _14336_/Q VGND VGND VPWR VPWR _13442_/X sky130_fd_sc_hd__mux2_1
X_10654_ _14757_/Q _10646_/X _10428_/X _10647_/X VGND VGND VPWR VPWR _14757_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13373_ _12634_/X _12611_/X _13418_/S VGND VGND VPWR VPWR _13373_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10585_ _10585_/A VGND VGND VPWR VPWR _10585_/X sky130_fd_sc_hd__buf_1
XFILLER_139_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15112_ _09270_/X _15112_/D VGND VGND VPWR VPWR _15112_/Q sky130_fd_sc_hd__dfxtp_1
X_12324_ _12324_/A _12324_/B VGND VGND VPWR VPWR _12325_/B sky130_fd_sc_hd__or2_1
XFILLER_5_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12255_ _12836_/A _12266_/B _12254_/Y VGND VGND VPWR VPWR _12798_/A sky130_fd_sc_hd__a21oi_1
X_15043_ _09518_/X _15043_/D VGND VGND VPWR VPWR _15043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11206_ _11219_/A VGND VGND VPWR VPWR _11207_/A sky130_fd_sc_hd__buf_1
X_12186_ _12190_/A VGND VGND VPWR VPWR _12762_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11137_ _11137_/A VGND VGND VPWR VPWR _11137_/X sky130_fd_sc_hd__clkbuf_1
X_11068_ _11068_/A VGND VGND VPWR VPWR _11068_/X sky130_fd_sc_hd__buf_1
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10019_ _10029_/A VGND VGND VPWR VPWR _10019_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14827_ _10402_/X _14827_/D VGND VGND VPWR VPWR _14827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14758_ _10651_/X _14758_/D VGND VGND VPWR VPWR _14758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13709_ _14845_/Q _14877_/Q _14909_/Q _14941_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13709_/X sky130_fd_sc_hd__mux4_2
XFILLER_149_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14689_ _10957_/X _14689_/D VGND VGND VPWR VPWR _14689_/Q sky130_fd_sc_hd__dfxtp_1
X_07230_ _07282_/B _07157_/B _07223_/X _07228_/Y VGND VGND VPWR VPWR _15643_/D sky130_fd_sc_hd__a211oi_2
XFILLER_20_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07161_ _07277_/B _07161_/B VGND VGND VPWR VPWR _07220_/A sky130_fd_sc_hd__or2_1
XFILLER_106_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09802_ _09802_/A VGND VGND VPWR VPWR _09802_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07994_ _07994_/A VGND VGND VPWR VPWR _07994_/X sky130_fd_sc_hd__buf_1
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09733_ _09733_/A VGND VGND VPWR VPWR _09754_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09664_ _15018_/Q _09660_/X _09662_/X _09663_/X VGND VGND VPWR VPWR _15018_/D sky130_fd_sc_hd__a22o_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08615_ _08635_/A VGND VGND VPWR VPWR _08622_/A sky130_fd_sc_hd__buf_1
XFILLER_43_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09595_ _10354_/A VGND VGND VPWR VPWR _09595_/X sky130_fd_sc_hd__buf_1
XFILLER_43_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08546_ _15299_/Q _08344_/A _08545_/X _08350_/A VGND VGND VPWR VPWR _15299_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08477_ _10775_/A VGND VGND VPWR VPWR _09245_/A sky130_fd_sc_hd__buf_1
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07428_ _07428_/A _13615_/X VGND VGND VPWR VPWR _15570_/D sky130_fd_sc_hd__and2_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07359_ _13153_/X _07298_/X _07498_/B _07354_/X _07358_/X VGND VGND VPWR VPWR _07362_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_149_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10370_ _10370_/A VGND VGND VPWR VPWR _10370_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09029_ _15174_/Q _09025_/X _08909_/X _09026_/X VGND VGND VPWR VPWR _15174_/D sky130_fd_sc_hd__a22o_1
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12040_ _12040_/A _12040_/B VGND VGND VPWR VPWR _12040_/X sky130_fd_sc_hd__or2_2
XFILLER_151_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13991_ _13987_/X _13988_/X _13989_/X _13990_/X _14397_/Q _14398_/Q VGND VGND VPWR
+ VPWR _13991_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12942_ _12692_/X _12703_/B _12957_/D _12938_/X _12941_/X VGND VGND VPWR VPWR _12942_/X
+ sky130_fd_sc_hd__o221a_1
X_15661_ _15663_/CLK _15661_/D VGND VGND VPWR VPWR _15661_/Q sky130_fd_sc_hd__dfxtp_1
X_12873_ _13314_/X VGND VGND VPWR VPWR _12873_/Y sky130_fd_sc_hd__inv_2
XANTENNA_110 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_121 rdata[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 rdata[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14612_ _11260_/X _14612_/D VGND VGND VPWR VPWR _14612_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_143 rdata[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11824_ _11828_/A VGND VGND VPWR VPWR _11824_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_154 rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15592_ _15592_/CLK _15592_/D VGND VGND VPWR VPWR _15592_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_165 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_176 wdata[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14543_ _11517_/X _14543_/D VGND VGND VPWR VPWR _14543_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_198 _13620_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11755_ _11755_/A VGND VGND VPWR VPWR _11820_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10706_ _10706_/A VGND VGND VPWR VPWR _10706_/X sky130_fd_sc_hd__clkbuf_1
X_14474_ _11773_/X _14474_/D VGND VGND VPWR VPWR _14474_/Q sky130_fd_sc_hd__dfxtp_1
X_11686_ _11686_/A _11798_/B VGND VGND VPWR VPWR _11700_/A sky130_fd_sc_hd__or2_2
XFILLER_146_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13425_ _12055_/Y _12983_/Y _13425_/S VGND VGND VPWR VPWR _13425_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10637_ _10646_/A VGND VGND VPWR VPWR _10637_/X sky130_fd_sc_hd__buf_1
XFILLER_139_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13356_ _12885_/X _12875_/B _13418_/S VGND VGND VPWR VPWR _13356_/X sky130_fd_sc_hd__mux2_1
X_10568_ _14783_/Q _10564_/X _10314_/X _10567_/X VGND VGND VPWR VPWR _14783_/D sky130_fd_sc_hd__a22o_1
XFILLER_115_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12307_ _12324_/A _12307_/B VGND VGND VPWR VPWR _12338_/A sky130_fd_sc_hd__or2_1
X_13287_ _13288_/X _13306_/X _15562_/Q VGND VGND VPWR VPWR _13287_/X sky130_fd_sc_hd__mux2_1
X_10499_ _10501_/A VGND VGND VPWR VPWR _10499_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15026_ _09615_/X _15026_/D VGND VGND VPWR VPWR _15026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12238_ _12238_/A VGND VGND VPWR VPWR _12239_/B sky130_fd_sc_hd__inv_2
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12169_ _12720_/A _12168_/A _12736_/A _12168_/Y VGND VGND VPWR VPWR _12685_/A sky130_fd_sc_hd__o22a_1
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08400_ _14327_/Q VGND VGND VPWR VPWR _10712_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09380_ _15084_/Q _09375_/X _09255_/X _09377_/X VGND VGND VPWR VPWR _15084_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08331_ _15334_/Q _08325_/X _08084_/X _08326_/X VGND VGND VPWR VPWR _15334_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08262_ _08262_/A VGND VGND VPWR VPWR _08262_/X sky130_fd_sc_hd__buf_1
X_07213_ _07268_/B _07167_/B _07212_/X _07208_/Y VGND VGND VPWR VPWR _15653_/D sky130_fd_sc_hd__a211oi_2
X_08193_ _08211_/A VGND VGND VPWR VPWR _08200_/A sky130_fd_sc_hd__buf_1
X_07144_ _13100_/X VGND VGND VPWR VPWR _07278_/B sky130_fd_sc_hd__inv_2
XFILLER_146_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07977_ _14327_/Q VGND VGND VPWR VPWR _07978_/A sky130_fd_sc_hd__buf_1
X_09716_ _09716_/A VGND VGND VPWR VPWR _09778_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_142_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09647_ _09647_/A VGND VGND VPWR VPWR _09647_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09578_ _10717_/A VGND VGND VPWR VPWR _10340_/A sky130_fd_sc_hd__buf_1
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _09279_/A VGND VGND VPWR VPWR _08529_/X sky130_fd_sc_hd__buf_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ _11552_/A VGND VGND VPWR VPWR _11540_/X sky130_fd_sc_hd__buf_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11471_ _11471_/A VGND VGND VPWR VPWR _11471_/X sky130_fd_sc_hd__buf_1
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ _13211_/X _13231_/X _15563_/Q VGND VGND VPWR VPWR _13210_/X sky130_fd_sc_hd__mux2_1
X_10422_ _10422_/A VGND VGND VPWR VPWR _10422_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14190_ _14957_/Q _15053_/Q _15021_/Q _15085_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14190_/X sky130_fd_sc_hd__mux4_2
XFILLER_136_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13141_ _12758_/A _13006_/Y _13152_/S VGND VGND VPWR VPWR _13141_/X sky130_fd_sc_hd__mux2_2
X_10353_ _10378_/A VGND VGND VPWR VPWR _10353_/X sky130_fd_sc_hd__buf_1
XFILLER_136_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13072_ _12732_/Y _15574_/Q _13076_/S VGND VGND VPWR VPWR _13072_/X sky130_fd_sc_hd__mux2_1
X_10284_ _10288_/A VGND VGND VPWR VPWR _10284_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12023_ _15513_/Q _12037_/A _15512_/Q _12023_/D VGND VGND VPWR VPWR _12024_/A sky130_fd_sc_hd__or4_4
XFILLER_78_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13974_ _15202_/Q _15170_/Q _14786_/Q _14818_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13974_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12925_ _12874_/Y _12879_/B _12869_/Y VGND VGND VPWR VPWR _12957_/C sky130_fd_sc_hd__o21ai_1
XFILLER_61_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15644_ _15646_/CLK _15644_/D VGND VGND VPWR VPWR _15644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12856_ _12699_/A _12854_/X _12829_/X _12855_/X VGND VGND VPWR VPWR _12856_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_61_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11807_ _11807_/A VGND VGND VPWR VPWR _11818_/A sky130_fd_sc_hd__clkbuf_2
X_15575_ _15576_/CLK _15575_/D VGND VGND VPWR VPWR _15575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12787_ _12745_/X _12777_/Y _12781_/Y _12786_/X VGND VGND VPWR VPWR _12787_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14526_ _11596_/X _14526_/D VGND VGND VPWR VPWR _14526_/Q sky130_fd_sc_hd__dfxtp_1
X_11738_ _11742_/A VGND VGND VPWR VPWR _11738_/X sky130_fd_sc_hd__clkbuf_1
X_14457_ _11833_/X _14457_/D VGND VGND VPWR VPWR _14457_/Q sky130_fd_sc_hd__dfxtp_1
X_11669_ _11669_/A VGND VGND VPWR VPWR _11669_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _13412_/X _13409_/X _13408_/S VGND VGND VPWR VPWR _13408_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14388_ _14399_/CLK instruction[25] VGND VGND VPWR VPWR _14388_/Q sky130_fd_sc_hd__dfxtp_4
X_13339_ _12875_/B _12885_/X _13418_/S VGND VGND VPWR VPWR _13339_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07900_ _07900_/A VGND VGND VPWR VPWR _07900_/Y sky130_fd_sc_hd__inv_2
X_15009_ _09707_/X _15009_/D VGND VGND VPWR VPWR _15009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08880_ _08906_/A VGND VGND VPWR VPWR _08880_/X sky130_fd_sc_hd__buf_1
X_07831_ _07872_/A _07831_/B _07831_/C VGND VGND VPWR VPWR _15449_/D sky130_fd_sc_hd__and3_1
XFILLER_57_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_opt_6_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR clkbuf_opt_6_clk/X sky130_fd_sc_hd__clkbuf_16
X_07762_ _07762_/A VGND VGND VPWR VPWR _07762_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09501_ _15049_/Q _09496_/X _09267_/X _09497_/X VGND VGND VPWR VPWR _15049_/D sky130_fd_sc_hd__a22o_1
X_07693_ _07652_/A _13129_/X _07652_/A _13129_/X VGND VGND VPWR VPWR _07827_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09432_ _15070_/Q _09425_/X _09176_/X _09428_/X VGND VGND VPWR VPWR _15070_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09363_ _09372_/A VGND VGND VPWR VPWR _09370_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08314_ _15339_/Q _08306_/X _08059_/X _08308_/X VGND VGND VPWR VPWR _15339_/D sky130_fd_sc_hd__a22o_1
X_09294_ _09923_/A _09294_/B _11574_/C VGND VGND VPWR VPWR _09810_/B sky130_fd_sc_hd__or3_1
XANTENNA_10 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08245_ _15359_/Q _08241_/X _07951_/X _08244_/X VGND VGND VPWR VPWR _15359_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_54 instruction[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_65 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_76 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08176_ _08178_/A VGND VGND VPWR VPWR _08176_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_98 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07127_ _13117_/X VGND VGND VPWR VPWR _07254_/B sky130_fd_sc_hd__inv_2
XFILLER_134_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10971_ _10975_/A VGND VGND VPWR VPWR _10971_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12710_ _12826_/A VGND VGND VPWR VPWR _12710_/X sky130_fd_sc_hd__buf_1
XFILLER_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13690_ _14975_/Q _15071_/Q _15039_/Q _15103_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13690_/X sky130_fd_sc_hd__mux4_2
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ _12641_/A _12641_/B VGND VGND VPWR VPWR _12641_/Y sky130_fd_sc_hd__nor2_1
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15360_ _08236_/X _15360_/D VGND VGND VPWR VPWR _15360_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12572_ _12572_/A _12572_/B VGND VGND VPWR VPWR _12572_/X sky130_fd_sc_hd__or2_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14311_ _14311_/CLK _14311_/D VGND VGND VPWR VPWR _14311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11523_ _11523_/A VGND VGND VPWR VPWR _11523_/X sky130_fd_sc_hd__buf_1
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15291_ _08579_/X _15291_/D VGND VGND VPWR VPWR _15291_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14242_ _15207_/Q _14535_/Q _14983_/Q _15399_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14242_/X sky130_fd_sc_hd__mux4_2
X_11454_ _11454_/A VGND VGND VPWR VPWR _11454_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10405_ _10410_/A VGND VGND VPWR VPWR _10405_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11385_ _11385_/A VGND VGND VPWR VPWR _11385_/X sky130_fd_sc_hd__buf_1
X_14173_ _14670_/Q _15246_/Q _14734_/Q _14702_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14173_/X sky130_fd_sc_hd__mux4_2
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13124_ _12435_/X _13023_/Y _13152_/S VGND VGND VPWR VPWR _13124_/X sky130_fd_sc_hd__mux2_2
X_10336_ _10336_/A VGND VGND VPWR VPWR _10336_/X sky130_fd_sc_hd__buf_1
XFILLER_3_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13055_ wdata[28] rdata[28] _13057_/S VGND VGND VPWR VPWR _14332_/D sky130_fd_sc_hd__mux2_1
X_10267_ _10280_/A VGND VGND VPWR VPWR _10267_/X sky130_fd_sc_hd__buf_1
XFILLER_79_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12006_ _12006_/A VGND VGND VPWR VPWR _12006_/X sky130_fd_sc_hd__buf_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10198_ _10258_/A VGND VGND VPWR VPWR _10218_/A sky130_fd_sc_hd__buf_2
XFILLER_78_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13957_ _14628_/Q _14596_/Q _14564_/Q _15364_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13957_/X sky130_fd_sc_hd__mux4_2
XFILLER_93_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12908_ _12908_/A _12908_/B _12949_/A _12908_/D VGND VGND VPWR VPWR _12909_/D sky130_fd_sc_hd__or4_4
XFILLER_74_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13888_ _14507_/Q _14475_/Q _14443_/Q _14411_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13888_/X sky130_fd_sc_hd__mux4_2
XFILLER_22_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15627_ _15669_/CLK _15627_/D VGND VGND VPWR VPWR pc[22] sky130_fd_sc_hd__dfxtp_4
XFILLER_22_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12839_ _12839_/A _12839_/B VGND VGND VPWR VPWR _12839_/Y sky130_fd_sc_hd__nand2_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15558_ _15589_/CLK _15558_/D VGND VGND VPWR VPWR _15558_/Q sky130_fd_sc_hd__dfxtp_1
X_14509_ _11650_/X _14509_/D VGND VGND VPWR VPWR _14509_/Q sky130_fd_sc_hd__dfxtp_1
X_15489_ _15510_/CLK _15489_/D VGND VGND VPWR VPWR wdata[15] sky130_fd_sc_hd__dfxtp_2
XFILLER_147_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08030_ _14317_/Q VGND VGND VPWR VPWR _08031_/A sky130_fd_sc_hd__buf_1
XFILLER_147_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09981_ _10349_/A VGND VGND VPWR VPWR _09981_/X sky130_fd_sc_hd__buf_1
XFILLER_131_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08932_ _08932_/A VGND VGND VPWR VPWR _08932_/X sky130_fd_sc_hd__buf_1
XFILLER_103_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08863_ _08868_/A VGND VGND VPWR VPWR _08863_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07814_ _07819_/A _07819_/B VGND VGND VPWR VPWR _07820_/B sky130_fd_sc_hd__or2_1
XFILLER_111_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08794_ _15232_/Q _08782_/X _08793_/X _08786_/X VGND VGND VPWR VPWR _15232_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07745_ _13147_/X VGND VGND VPWR VPWR _07746_/A sky130_fd_sc_hd__inv_2
XFILLER_84_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07676_ _07781_/A _07674_/X _07675_/X _13128_/X VGND VGND VPWR VPWR _07819_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09415_ _09508_/A VGND VGND VPWR VPWR _09478_/A sky130_fd_sc_hd__buf_1
XFILLER_25_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09346_ _09376_/A VGND VGND VPWR VPWR _09366_/A sky130_fd_sc_hd__buf_2
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09277_ _15111_/Q _09274_/X _09275_/X _09276_/X VGND VGND VPWR VPWR _15111_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08228_ _08239_/A VGND VGND VPWR VPWR _08242_/A sky130_fd_sc_hd__inv_2
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08159_ _08159_/A VGND VGND VPWR VPWR _08159_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11170_ _11537_/A VGND VGND VPWR VPWR _11170_/X sky130_fd_sc_hd__buf_1
X_10121_ _10123_/A VGND VGND VPWR VPWR _10121_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10052_ _10052_/A VGND VGND VPWR VPWR _10052_/X sky130_fd_sc_hd__buf_1
XFILLER_0_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14860_ _10262_/X _14860_/D VGND VGND VPWR VPWR _14860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13811_ _13807_/X _13808_/X _13809_/X _13810_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13811_/X sky130_fd_sc_hd__mux4_2
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14791_ _10534_/X _14791_/D VGND VGND VPWR VPWR _14791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13742_ _15225_/Q _14553_/Q _15001_/Q _15417_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13742_/X sky130_fd_sc_hd__mux4_1
X_10954_ _10954_/A VGND VGND VPWR VPWR _10954_/X sky130_fd_sc_hd__buf_1
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13673_ _14688_/Q _15264_/Q _14752_/Q _14720_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13673_/X sky130_fd_sc_hd__mux4_2
X_10885_ _10915_/A VGND VGND VPWR VPWR _10905_/A sky130_fd_sc_hd__buf_1
XFILLER_31_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15412_ _08009_/X _15412_/D VGND VGND VPWR VPWR _15412_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12624_ _12578_/X _12614_/Y _12617_/Y _12619_/X _12623_/X VGND VGND VPWR VPWR _12624_/Y
+ sky130_fd_sc_hd__o2111ai_4
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15343_ _08300_/X _15343_/D VGND VGND VPWR VPWR _15343_/Q sky130_fd_sc_hd__dfxtp_1
X_12555_ _15471_/Q _12550_/Y data_address[0] VGND VGND VPWR VPWR _12561_/B sky130_fd_sc_hd__a21oi_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11506_ _11506_/A VGND VGND VPWR VPWR _11506_/X sky130_fd_sc_hd__buf_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15274_ _08636_/X _15274_/D VGND VGND VPWR VPWR _15274_/Q sky130_fd_sc_hd__dfxtp_1
X_12486_ _12519_/A VGND VGND VPWR VPWR _12796_/A sky130_fd_sc_hd__clkbuf_2
X_14225_ _15113_/Q _15337_/Q _15305_/Q _15273_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14225_/X sky130_fd_sc_hd__mux4_1
X_11437_ _11437_/A VGND VGND VPWR VPWR _11437_/X sky130_fd_sc_hd__buf_1
XFILLER_125_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14156_ _14152_/X _14153_/X _14154_/X _14155_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14156_/X sky130_fd_sc_hd__mux4_2
X_11368_ _11368_/A VGND VGND VPWR VPWR _11373_/A sky130_fd_sc_hd__buf_2
XFILLER_98_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13107_ _15653_/Q data_address[18] _15667_/Q VGND VGND VPWR VPWR _13107_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10319_ _10319_/A VGND VGND VPWR VPWR _10319_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14087_ _14647_/Q _14615_/Q _14583_/Q _15383_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14087_/X sky130_fd_sc_hd__mux4_2
X_11299_ _11299_/A VGND VGND VPWR VPWR _11299_/X sky130_fd_sc_hd__clkbuf_1
X_13038_ wdata[11] rdata[11] ren VGND VGND VPWR VPWR _14315_/D sky130_fd_sc_hd__mux2_2
XFILLER_39_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14989_ _09775_/X _14989_/D VGND VGND VPWR VPWR _14989_/Q sky130_fd_sc_hd__dfxtp_1
X_07530_ _15470_/Q VGND VGND VPWR VPWR _07530_/Y sky130_fd_sc_hd__inv_2
X_07461_ _07469_/A VGND VGND VPWR VPWR _07464_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_90_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09200_ _09200_/A VGND VGND VPWR VPWR _09200_/X sky130_fd_sc_hd__buf_1
XFILLER_50_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07392_ _07491_/A _07392_/B VGND VGND VPWR VPWR _15593_/D sky130_fd_sc_hd__nor2_1
XFILLER_22_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09131_ _09135_/A VGND VGND VPWR VPWR _09131_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09062_ _09064_/A VGND VGND VPWR VPWR _09062_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08013_ _08019_/A VGND VGND VPWR VPWR _08013_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09964_ _09964_/A VGND VGND VPWR VPWR _10173_/A sky130_fd_sc_hd__buf_1
XFILLER_89_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08915_ _08918_/A VGND VGND VPWR VPWR _08915_/X sky130_fd_sc_hd__clkbuf_1
X_09895_ _09897_/A VGND VGND VPWR VPWR _09895_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08846_ _08846_/A VGND VGND VPWR VPWR _08855_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08777_ _08788_/A VGND VGND VPWR VPWR _08777_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07728_ _13143_/X _07728_/B VGND VGND VPWR VPWR _07728_/Y sky130_fd_sc_hd__nor2_1
X_07659_ _07848_/A VGND VGND VPWR VPWR _07659_/X sky130_fd_sc_hd__buf_1
XFILLER_40_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10670_ _10670_/A VGND VGND VPWR VPWR _10670_/X sky130_fd_sc_hd__clkbuf_1
X_09329_ _09331_/A VGND VGND VPWR VPWR _09329_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12340_ _12417_/A VGND VGND VPWR VPWR _12493_/A sky130_fd_sc_hd__buf_1
XFILLER_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12271_ _12271_/A _12271_/B VGND VGND VPWR VPWR _12271_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14010_ _14975_/Q _15071_/Q _15039_/Q _15103_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14010_/X sky130_fd_sc_hd__mux4_2
X_11222_ _11222_/A VGND VGND VPWR VPWR _11285_/A sky130_fd_sc_hd__buf_2
XFILLER_108_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11153_ _14639_/Q _11147_/X _11152_/X _11149_/X VGND VGND VPWR VPWR _14639_/D sky130_fd_sc_hd__a22o_1
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10104_ _10104_/A VGND VGND VPWR VPWR _10111_/A sky130_fd_sc_hd__buf_1
X_11084_ _11109_/A VGND VGND VPWR VPWR _11084_/X sky130_fd_sc_hd__buf_1
XFILLER_150_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14912_ _10078_/X _14912_/D VGND VGND VPWR VPWR _14912_/Q sky130_fd_sc_hd__dfxtp_1
X_10035_ _14923_/Q _10024_/X _10034_/X _10027_/X VGND VGND VPWR VPWR _14923_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14843_ _10331_/X _14843_/D VGND VGND VPWR VPWR _14843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14774_ _10595_/X _14774_/D VGND VGND VPWR VPWR _14774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11986_ _12005_/A VGND VGND VPWR VPWR _11986_/X sky130_fd_sc_hd__buf_1
XFILLER_91_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13725_ _15131_/Q _15355_/Q _15323_/Q _15291_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13725_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10937_ _10937_/A VGND VGND VPWR VPWR _10937_/X sky130_fd_sc_hd__buf_1
XFILLER_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13656_ _13652_/X _13653_/X _13654_/X _13655_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13656_/X sky130_fd_sc_hd__mux4_2
X_10868_ _14715_/Q _10864_/X _10708_/X _10865_/X VGND VGND VPWR VPWR _14715_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12607_ _12371_/A _12604_/Y _13204_/X _12417_/A _12606_/Y VGND VGND VPWR VPWR _12607_/X
+ sky130_fd_sc_hd__o221a_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13587_ _13586_/X _13075_/X _14337_/Q VGND VGND VPWR VPWR _13587_/X sky130_fd_sc_hd__mux2_1
X_10799_ _11541_/A VGND VGND VPWR VPWR _10799_/X sky130_fd_sc_hd__buf_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15326_ _08374_/X _15326_/D VGND VGND VPWR VPWR _15326_/Q sky130_fd_sc_hd__dfxtp_1
X_12538_ _15462_/Q _15461_/Q _15463_/Q _15465_/Q VGND VGND VPWR VPWR _12538_/X sky130_fd_sc_hd__or4_4
XFILLER_8_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15257_ _08701_/X _15257_/D VGND VGND VPWR VPWR _15257_/Q sky130_fd_sc_hd__dfxtp_1
X_12469_ _12467_/Y _12468_/X _12467_/Y _12468_/X VGND VGND VPWR VPWR _12469_/Y sky130_fd_sc_hd__a2bb2oi_2
X_14208_ _14507_/Q _14475_/Q _14443_/Q _14411_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14208_/X sky130_fd_sc_hd__mux4_2
XFILLER_126_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15188_ _08980_/X _15188_/D VGND VGND VPWR VPWR _15188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14139_ _14834_/Q _14866_/Q _14898_/Q _14930_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14139_/X sky130_fd_sc_hd__mux4_2
XFILLER_113_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08700_ _15258_/Q _08693_/X _08402_/X _08694_/X VGND VGND VPWR VPWR _15258_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09680_ _09680_/A VGND VGND VPWR VPWR _09680_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08631_ _08633_/A VGND VGND VPWR VPWR _08631_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08562_ _08572_/A VGND VGND VPWR VPWR _08562_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07513_ _07514_/A _07513_/B VGND VGND VPWR VPWR _15513_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08493_ _15308_/Q _08482_/X _08492_/X _08487_/X VGND VGND VPWR VPWR _15308_/D sky130_fd_sc_hd__a22o_1
X_07444_ _07446_/A _13430_/X VGND VGND VPWR VPWR _15560_/D sky130_fd_sc_hd__and2_1
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07375_ _13155_/X _07363_/X _07508_/B _07354_/X _07374_/X VGND VGND VPWR VPWR _07377_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_50_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09114_ _09114_/A VGND VGND VPWR VPWR _09114_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09045_ _15170_/Q _09041_/X _08783_/X _09044_/X VGND VGND VPWR VPWR _15170_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09947_ _09974_/A VGND VGND VPWR VPWR _09947_/X sky130_fd_sc_hd__buf_1
XFILLER_131_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09878_ _09878_/A VGND VGND VPWR VPWR _09878_/X sky130_fd_sc_hd__buf_1
XFILLER_100_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08829_ _08829_/A VGND VGND VPWR VPWR _08829_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11840_ _11848_/A VGND VGND VPWR VPWR _11840_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11771_ _11773_/A VGND VGND VPWR VPWR _11771_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13510_ _13509_/X rdata[4] _14338_/Q VGND VGND VPWR VPWR _13510_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10722_ _10722_/A VGND VGND VPWR VPWR _11479_/A sky130_fd_sc_hd__buf_1
X_14490_ _11719_/X _14490_/D VGND VGND VPWR VPWR _14490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13441_ _13440_/X rdata[27] _13516_/S VGND VGND VPWR VPWR _13441_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10653_ _10655_/A VGND VGND VPWR VPWR _10653_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13372_ _13374_/X _13373_/X _13415_/S VGND VGND VPWR VPWR _13372_/X sky130_fd_sc_hd__mux2_1
X_10584_ _10584_/A VGND VGND VPWR VPWR _10584_/X sky130_fd_sc_hd__buf_1
X_15111_ _09273_/X _15111_/D VGND VGND VPWR VPWR _15111_/Q sky130_fd_sc_hd__dfxtp_1
X_12323_ _12878_/A _13394_/X VGND VGND VPWR VPWR _12323_/X sky130_fd_sc_hd__or2_2
XFILLER_5_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15042_ _09520_/X _15042_/D VGND VGND VPWR VPWR _15042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12254_ _12254_/A _12266_/B VGND VGND VPWR VPWR _12254_/Y sky130_fd_sc_hd__nor2_1
X_11205_ _11317_/A _11428_/B VGND VGND VPWR VPWR _11219_/A sky130_fd_sc_hd__or2_2
XFILLER_135_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12185_ _15539_/Q VGND VGND VPWR VPWR _12190_/A sky130_fd_sc_hd__inv_2
X_11136_ _14643_/Q _11133_/X _11134_/X _11135_/X VGND VGND VPWR VPWR _14643_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11067_ _11082_/A VGND VGND VPWR VPWR _11068_/A sky130_fd_sc_hd__buf_1
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10018_ _10032_/A VGND VGND VPWR VPWR _10029_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14826_ _10405_/X _14826_/D VGND VGND VPWR VPWR _14826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14757_ _10653_/X _14757_/D VGND VGND VPWR VPWR _14757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11969_ _11971_/A VGND VGND VPWR VPWR _11969_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13708_ _14525_/Q _14493_/Q _14461_/Q _14429_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13708_/X sky130_fd_sc_hd__mux4_2
XFILLER_60_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14688_ _10959_/X _14688_/D VGND VGND VPWR VPWR _14688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13639_ _13638_/X _13062_/X _14337_/Q VGND VGND VPWR VPWR _13639_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07160_ _07278_/B _07225_/A VGND VGND VPWR VPWR _07161_/B sky130_fd_sc_hd__or2_1
XFILLER_145_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15309_ _08480_/X _15309_/D VGND VGND VPWR VPWR _15309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09801_ _14982_/Q _09797_/X _09682_/X _09798_/X VGND VGND VPWR VPWR _14982_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07993_ _14324_/Q VGND VGND VPWR VPWR _07994_/A sky130_fd_sc_hd__buf_1
XFILLER_101_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09732_ _15002_/Q _09726_/X _09574_/X _09727_/X VGND VGND VPWR VPWR _15002_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09663_ _09678_/A VGND VGND VPWR VPWR _09663_/X sky130_fd_sc_hd__buf_1
XFILLER_28_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08614_ _08644_/A VGND VGND VPWR VPWR _08635_/A sky130_fd_sc_hd__buf_4
XFILLER_43_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09594_ _10733_/A VGND VGND VPWR VPWR _10354_/A sky130_fd_sc_hd__buf_1
XFILLER_82_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08545_ _09290_/A VGND VGND VPWR VPWR _08545_/X sky130_fd_sc_hd__buf_1
XFILLER_70_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08476_ _14315_/Q VGND VGND VPWR VPWR _10775_/A sky130_fd_sc_hd__buf_1
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07427_ _07428_/A _13611_/X VGND VGND VPWR VPWR _15571_/D sky130_fd_sc_hd__and2_1
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07358_ _07506_/B _07356_/X _12574_/A _07308_/X VGND VGND VPWR VPWR _07358_/X sky130_fd_sc_hd__o22a_1
X_07289_ _15637_/D VGND VGND VPWR VPWR _15607_/D sky130_fd_sc_hd__inv_2
XFILLER_108_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09028_ _09030_/A VGND VGND VPWR VPWR _09028_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13990_ _14977_/Q _15073_/Q _15041_/Q _15105_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13990_/X sky130_fd_sc_hd__mux4_2
XFILLER_86_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12941_ _12941_/A _12941_/B VGND VGND VPWR VPWR _12941_/X sky130_fd_sc_hd__or2_1
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15660_ _15663_/CLK _15660_/D VGND VGND VPWR VPWR _15660_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_100 pc[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12872_ _12707_/A _12861_/X _12663_/X _12865_/Y _12871_/X VGND VGND VPWR VPWR _12872_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA_111 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14611_ _11263_/X _14611_/D VGND VGND VPWR VPWR _14611_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_122 rdata[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_133 rdata[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11823_ _14461_/Q _11813_/X _07963_/A _11816_/X VGND VGND VPWR VPWR _14461_/D sky130_fd_sc_hd__a22o_1
XANTENNA_144 rdata[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15591_ _15591_/CLK _15591_/D VGND VGND VPWR VPWR _15591_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_155 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14542_ _11522_/X _14542_/D VGND VGND VPWR VPWR _14542_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_177 wdata[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11754_ _14480_/Q _11752_/X _11514_/X _11753_/X VGND VGND VPWR VPWR _14480_/D sky130_fd_sc_hd__a22o_1
XANTENNA_188 wdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_199 _13616_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10705_ _14748_/Q _10701_/X _10703_/X _10704_/X VGND VGND VPWR VPWR _14748_/D sky130_fd_sc_hd__a22o_1
X_14473_ _11778_/X _14473_/D VGND VGND VPWR VPWR _14473_/Q sky130_fd_sc_hd__dfxtp_1
X_11685_ _11685_/A VGND VGND VPWR VPWR _11685_/X sky130_fd_sc_hd__clkbuf_1
X_13424_ _15520_/Q _15521_/Q _15519_/Q VGND VGND VPWR VPWR _13424_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10636_ _10636_/A VGND VGND VPWR VPWR _10636_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13355_ _12885_/X _12817_/B _15561_/Q VGND VGND VPWR VPWR _13355_/X sky130_fd_sc_hd__mux2_1
X_10567_ _10585_/A VGND VGND VPWR VPWR _10567_/X sky130_fd_sc_hd__buf_1
XFILLER_6_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12306_ _12316_/B _12324_/B VGND VGND VPWR VPWR _12333_/A sky130_fd_sc_hd__or2_1
XFILLER_127_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13286_ _13287_/X _13322_/X _15563_/Q VGND VGND VPWR VPWR _13286_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10498_ _14803_/Q _10496_/X _10367_/X _10497_/X VGND VGND VPWR VPWR _14803_/D sky130_fd_sc_hd__a22o_1
X_15025_ _09620_/X _15025_/D VGND VGND VPWR VPWR _15025_/Q sky130_fd_sc_hd__dfxtp_1
X_12237_ _12235_/X _12157_/A _12807_/A _12105_/A VGND VGND VPWR VPWR _12238_/A sky130_fd_sc_hd__o22a_1
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12168_ _12168_/A VGND VGND VPWR VPWR _12168_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11119_ _11159_/A VGND VGND VPWR VPWR _11147_/A sky130_fd_sc_hd__buf_2
X_12099_ _15550_/Q VGND VGND VPWR VPWR _12109_/A sky130_fd_sc_hd__inv_2
XFILLER_96_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14809_ _10473_/X _14809_/D VGND VGND VPWR VPWR _14809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08330_ _08334_/A VGND VGND VPWR VPWR _08330_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08261_ _08261_/A VGND VGND VPWR VPWR _08261_/X sky130_fd_sc_hd__buf_1
XFILLER_119_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07212_ _07246_/A VGND VGND VPWR VPWR _07212_/X sky130_fd_sc_hd__buf_2
X_08192_ _08264_/A VGND VGND VPWR VPWR _08211_/A sky130_fd_sc_hd__buf_1
X_07143_ _13101_/X VGND VGND VPWR VPWR _07277_/B sky130_fd_sc_hd__inv_2
XFILLER_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07976_ _07986_/A VGND VGND VPWR VPWR _07976_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09715_ _09736_/A VGND VGND VPWR VPWR _09715_/X sky130_fd_sc_hd__buf_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09646_ _15021_/Q _09641_/X _09643_/X _09645_/X VGND VGND VPWR VPWR _15021_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09577_ _09577_/A VGND VGND VPWR VPWR _09577_/X sky130_fd_sc_hd__buf_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08528_ _10818_/A VGND VGND VPWR VPWR _09279_/A sky130_fd_sc_hd__buf_1
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _10760_/A VGND VGND VPWR VPWR _09232_/A sky130_fd_sc_hd__clkbuf_2
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ _11478_/A VGND VGND VPWR VPWR _11470_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10421_ _14823_/Q _10418_/X _10419_/X _10420_/X VGND VGND VPWR VPWR _14823_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13140_ _12737_/A _13007_/Y _13152_/S VGND VGND VPWR VPWR _13140_/X sky130_fd_sc_hd__mux2_1
X_10352_ _10392_/A VGND VGND VPWR VPWR _10378_/A sky130_fd_sc_hd__buf_2
XFILLER_109_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13071_ _12744_/X _15573_/Q _13076_/S VGND VGND VPWR VPWR _13071_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10283_ _10290_/A VGND VGND VPWR VPWR _10288_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12022_ _15511_/Q VGND VGND VPWR VPWR _12037_/A sky130_fd_sc_hd__inv_2
XFILLER_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13973_ _14690_/Q _15266_/Q _14754_/Q _14722_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _13973_/X sky130_fd_sc_hd__mux4_2
XFILLER_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12924_ _12924_/A _12924_/B _12924_/C _12933_/A VGND VGND VPWR VPWR _12958_/B sky130_fd_sc_hd__or4_4
XFILLER_46_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12855_ _12852_/X _12838_/X _12830_/X VGND VGND VPWR VPWR _12855_/X sky130_fd_sc_hd__o21a_1
X_15643_ _15647_/CLK _15643_/D VGND VGND VPWR VPWR _15643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11806_ _14465_/Q _11800_/X _07936_/A _11803_/X VGND VGND VPWR VPWR _14465_/D sky130_fd_sc_hd__a22o_1
X_15574_ _15576_/CLK _15574_/D VGND VGND VPWR VPWR _15574_/Q sky130_fd_sc_hd__dfxtp_1
X_12786_ _13279_/X _12782_/X _13274_/X _12810_/A _12785_/X VGND VGND VPWR VPWR _12786_/X
+ sky130_fd_sc_hd__o221a_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14525_ _11598_/X _14525_/D VGND VGND VPWR VPWR _14525_/Q sky130_fd_sc_hd__dfxtp_1
X_11737_ _11746_/A VGND VGND VPWR VPWR _11742_/A sky130_fd_sc_hd__buf_1
XFILLER_30_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14456_ _11837_/X _14456_/D VGND VGND VPWR VPWR _14456_/Q sky130_fd_sc_hd__dfxtp_1
X_11668_ _14505_/Q _11664_/X _11545_/X _11665_/X VGND VGND VPWR VPWR _14505_/D sky130_fd_sc_hd__a22o_1
XFILLER_128_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _12662_/X _12138_/X _13418_/S VGND VGND VPWR VPWR _13407_/X sky130_fd_sc_hd__mux2_1
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10619_ _10649_/A VGND VGND VPWR VPWR _10640_/A sky130_fd_sc_hd__clkbuf_2
X_14387_ _14395_/CLK instruction[24] VGND VGND VPWR VPWR _14387_/Q sky130_fd_sc_hd__dfxtp_4
X_11599_ _14525_/Q _11591_/X _11459_/X _11594_/X VGND VGND VPWR VPWR _14525_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13338_ _12882_/Y _12926_/B _13415_/S VGND VGND VPWR VPWR _13338_/X sky130_fd_sc_hd__mux2_1
X_13269_ _13270_/X _13296_/X _13408_/S VGND VGND VPWR VPWR _13269_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15008_ _09709_/X _15008_/D VGND VGND VPWR VPWR _15008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07830_ _07830_/A _07830_/B VGND VGND VPWR VPWR _07831_/C sky130_fd_sc_hd__nand2_1
XFILLER_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07761_ _13151_/X _07757_/Y _07909_/B VGND VGND VPWR VPWR _07762_/A sky130_fd_sc_hd__o21ai_2
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09500_ _09504_/A VGND VGND VPWR VPWR _09500_/X sky130_fd_sc_hd__clkbuf_1
X_07692_ _07689_/X _07688_/X _07689_/X _13130_/X VGND VGND VPWR VPWR _07830_/A sky130_fd_sc_hd__a2bb2o_1
X_09431_ _09435_/A VGND VGND VPWR VPWR _09431_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09362_ _15089_/Q _09356_/X _09232_/X _09357_/X VGND VGND VPWR VPWR _15089_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08313_ _08315_/A VGND VGND VPWR VPWR _08313_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09293_ _09305_/A VGND VGND VPWR VPWR _09293_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_11 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_22 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_33 data_address[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08244_ _08262_/A VGND VGND VPWR VPWR _08244_/X sky130_fd_sc_hd__buf_1
XANTENNA_44 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 instruction[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_66 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08175_ _15376_/Q _08173_/X _08031_/X _08174_/X VGND VGND VPWR VPWR _15376_/D sky130_fd_sc_hd__a22o_1
XANTENNA_88 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_99 pc[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07126_ _13118_/X VGND VGND VPWR VPWR _07252_/B sky130_fd_sc_hd__inv_2
XFILLER_134_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07959_ _15422_/Q _07949_/X _07958_/X _07954_/X VGND VGND VPWR VPWR _15422_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10970_ _10988_/A VGND VGND VPWR VPWR _10975_/A sky130_fd_sc_hd__buf_1
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09629_ _15024_/Q _09625_/X _09627_/X _09628_/X VGND VGND VPWR VPWR _15024_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ _12640_/A VGND VGND VPWR VPWR _12640_/Y sky130_fd_sc_hd__inv_2
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12571_ _12571_/A VGND VGND VPWR VPWR _12572_/A sky130_fd_sc_hd__buf_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_50_clk _14315_/CLK VGND VGND VPWR VPWR _15666_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ _14311_/CLK _14310_/D VGND VGND VPWR VPWR _14310_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ _11532_/A VGND VGND VPWR VPWR _11522_/X sky130_fd_sc_hd__clkbuf_2
X_15290_ _08581_/X _15290_/D VGND VGND VPWR VPWR _15290_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14241_ _14237_/X _14238_/X _14239_/X _14240_/X _14266_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14241_/X sky130_fd_sc_hd__mux4_1
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11453_ _14559_/Q _11448_/X _11449_/X _11452_/X VGND VGND VPWR VPWR _14559_/D sky130_fd_sc_hd__a22o_1
X_10404_ _14827_/Q _10393_/X _10403_/X _10396_/X VGND VGND VPWR VPWR _14827_/D sky130_fd_sc_hd__a22o_1
X_14172_ _15214_/Q _14542_/Q _14990_/Q _15406_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14172_/X sky130_fd_sc_hd__mux4_2
X_11384_ _11384_/A VGND VGND VPWR VPWR _11384_/X sky130_fd_sc_hd__buf_1
XFILLER_109_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13123_ _12480_/B _13024_/Y _13152_/S VGND VGND VPWR VPWR _13123_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10335_ _10343_/A VGND VGND VPWR VPWR _10335_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13054_ wdata[27] rdata[27] _13057_/S VGND VGND VPWR VPWR _14331_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10266_ _10266_/A VGND VGND VPWR VPWR _10266_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12005_ _12005_/A VGND VGND VPWR VPWR _12005_/X sky130_fd_sc_hd__buf_1
XFILLER_78_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10197_ _10197_/A VGND VGND VPWR VPWR _10258_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13956_ _13952_/X _13953_/X _13954_/X _13955_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13956_/X sky130_fd_sc_hd__mux4_2
X_12907_ _12132_/X _15577_/Q _12661_/A _12676_/A VGND VGND VPWR VPWR _12908_/D sky130_fd_sc_hd__o22a_1
XFILLER_61_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13887_ _14635_/Q _14603_/Q _14571_/Q _15371_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13887_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12838_ _12838_/A VGND VGND VPWR VPWR _12838_/X sky130_fd_sc_hd__clkbuf_4
X_15626_ _15662_/CLK _15626_/D VGND VGND VPWR VPWR pc[21] sky130_fd_sc_hd__dfxtp_4
XFILLER_62_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12769_ _13268_/X _12707_/X _12764_/X _12767_/Y _12768_/Y VGND VGND VPWR VPWR _12769_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_15_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15557_ _15589_/CLK _15557_/D VGND VGND VPWR VPWR _15557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR _15517_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14508_ _11656_/X _14508_/D VGND VGND VPWR VPWR _14508_/Q sky130_fd_sc_hd__dfxtp_1
X_15488_ _15667_/CLK _15488_/D VGND VGND VPWR VPWR wdata[14] sky130_fd_sc_hd__dfxtp_2
X_14439_ _11894_/X _14439_/D VGND VGND VPWR VPWR _14439_/Q sky130_fd_sc_hd__dfxtp_1
X_09980_ _09990_/A VGND VGND VPWR VPWR _09980_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08931_ _08944_/A VGND VGND VPWR VPWR _08932_/A sky130_fd_sc_hd__buf_1
XFILLER_130_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08862_ _15217_/Q _08851_/X _08861_/X _08853_/X VGND VGND VPWR VPWR _15217_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07813_ _07848_/A VGND VGND VPWR VPWR _07813_/X sky130_fd_sc_hd__buf_1
X_08793_ _09164_/A VGND VGND VPWR VPWR _08793_/X sky130_fd_sc_hd__buf_1
XFILLER_38_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07744_ _13146_/X _07742_/Y _07743_/Y _15599_/Q VGND VGND VPWR VPWR _07889_/B sky130_fd_sc_hd__o22a_1
XFILLER_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07675_ _07675_/A VGND VGND VPWR VPWR _07675_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09414_ _15074_/Q _09410_/X _09153_/X _09413_/X VGND VGND VPWR VPWR _15074_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09345_ _09365_/A VGND VGND VPWR VPWR _09345_/X sky130_fd_sc_hd__buf_1
XFILLER_40_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk _14315_/CLK VGND VGND VPWR VPWR _15646_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09276_ _09276_/A VGND VGND VPWR VPWR _09276_/X sky130_fd_sc_hd__buf_1
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08227_ _08227_/A VGND VGND VPWR VPWR _08227_/X sky130_fd_sc_hd__buf_1
XFILLER_138_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08158_ _15381_/Q _08153_/X _08006_/X _08155_/X VGND VGND VPWR VPWR _15381_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07109_ _07795_/A VGND VGND VPWR VPWR _07893_/A sky130_fd_sc_hd__buf_1
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08089_ _08097_/A VGND VGND VPWR VPWR _08089_/X sky130_fd_sc_hd__buf_1
XFILLER_134_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10120_ _14902_/Q _10117_/X _09986_/X _10119_/X VGND VGND VPWR VPWR _14902_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10051_ _10419_/A VGND VGND VPWR VPWR _10051_/X sky130_fd_sc_hd__buf_1
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13810_ _14963_/Q _15059_/Q _15027_/Q _15091_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13810_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14790_ _10538_/X _14790_/D VGND VGND VPWR VPWR _14790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13741_ _13737_/X _13738_/X _13739_/X _13740_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13741_/X sky130_fd_sc_hd__mux4_1
X_10953_ _10965_/A VGND VGND VPWR VPWR _10954_/A sky130_fd_sc_hd__buf_1
XFILLER_44_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13672_ _15232_/Q _14560_/Q _15008_/Q _15424_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13672_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10884_ _10904_/A VGND VGND VPWR VPWR _10884_/X sky130_fd_sc_hd__buf_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15411_ _08013_/X _15411_/D VGND VGND VPWR VPWR _15411_/Q sky130_fd_sc_hd__dfxtp_1
X_12623_ _13310_/X _12620_/X _12593_/X _12622_/Y VGND VGND VPWR VPWR _12623_/X sky130_fd_sc_hd__o22a_1
XFILLER_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_clk _14328_/CLK VGND VGND VPWR VPWR _15589_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15342_ _08302_/X _15342_/D VGND VGND VPWR VPWR _15342_/Q sky130_fd_sc_hd__dfxtp_1
X_12554_ _12546_/X _12549_/Y _12553_/X VGND VGND VPWR VPWR wstrobe[0] sky130_fd_sc_hd__o21a_2
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11505_ _11505_/A VGND VGND VPWR VPWR _11505_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15273_ _08640_/X _15273_/D VGND VGND VPWR VPWR _15273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12485_ _15562_/Q VGND VGND VPWR VPWR _12519_/A sky130_fd_sc_hd__buf_1
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14224_ _15177_/Q _15145_/Q _14761_/Q _14793_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14224_/X sky130_fd_sc_hd__mux4_2
XFILLER_144_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11436_ _11436_/A VGND VGND VPWR VPWR _11436_/X sky130_fd_sc_hd__clkbuf_1
X_14155_ _15120_/Q _15344_/Q _15312_/Q _15280_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14155_/X sky130_fd_sc_hd__mux4_2
X_11367_ _14582_/Q _11364_/X _11121_/X _11366_/X VGND VGND VPWR VPWR _14582_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13106_ _15652_/Q data_address[17] _15667_/Q VGND VGND VPWR VPWR _13106_/X sky130_fd_sc_hd__mux2_1
X_10318_ _14847_/Q _10313_/X _10314_/X _10317_/X VGND VGND VPWR VPWR _14847_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14086_ _14082_/X _14083_/X _14084_/X _14085_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14086_/X sky130_fd_sc_hd__mux4_2
X_11298_ _14601_/Q _11294_/X _11178_/X _11295_/X VGND VGND VPWR VPWR _14601_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13037_ wdata[10] rdata[10] ren VGND VGND VPWR VPWR _14314_/D sky130_fd_sc_hd__mux2_4
XFILLER_79_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10249_ _14864_/Q _10247_/X _10012_/X _10248_/X VGND VGND VPWR VPWR _14864_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14988_ _09781_/X _14988_/D VGND VGND VPWR VPWR _14988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13939_ _14822_/Q _14854_/Q _14886_/Q _14918_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13939_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07460_ _07460_/A VGND VGND VPWR VPWR _07469_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15609_ _15648_/CLK _15609_/D VGND VGND VPWR VPWR pc[4] sky130_fd_sc_hd__dfxtp_1
X_07391_ _07392_/B VGND VGND VPWR VPWR _07391_/Y sky130_fd_sc_hd__inv_2
X_09130_ _09146_/A VGND VGND VPWR VPWR _09135_/A sky130_fd_sc_hd__buf_1
XFILLER_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09061_ _15166_/Q _09054_/X _08805_/X _09057_/X VGND VGND VPWR VPWR _15166_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08012_ _15412_/Q _07998_/X _08011_/X _08002_/X VGND VGND VPWR VPWR _15412_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09963_ _14939_/Q _09957_/X _09962_/X _09959_/X VGND VGND VPWR VPWR _14939_/D sky130_fd_sc_hd__a22o_1
X_08914_ _15205_/Q _08904_/X _08913_/X _08906_/X VGND VGND VPWR VPWR _15205_/D sky130_fd_sc_hd__a22o_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09894_ _14956_/Q _09887_/X _09649_/X _09889_/X VGND VGND VPWR VPWR _14956_/D sky130_fd_sc_hd__a22o_1
XFILLER_131_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08845_ _15221_/Q _08838_/X _08844_/X _08841_/X VGND VGND VPWR VPWR _15221_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08776_ _15235_/Q _08666_/A _08545_/X _08669_/A VGND VGND VPWR VPWR _15235_/D sky130_fd_sc_hd__a22o_1
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07727_ _15602_/Q VGND VGND VPWR VPWR _07728_/B sky130_fd_sc_hd__inv_2
XFILLER_81_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07658_ _07658_/A VGND VGND VPWR VPWR _07848_/A sky130_fd_sc_hd__buf_1
XFILLER_26_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07589_ _07591_/A _13076_/X VGND VGND VPWR VPWR _15491_/D sky130_fd_sc_hd__and2_1
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09328_ _15100_/Q _09326_/X _09184_/X _09327_/X VGND VGND VPWR VPWR _15100_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09259_ _09259_/A VGND VGND VPWR VPWR _09259_/X sky130_fd_sc_hd__buf_1
XFILLER_139_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12270_ _12800_/A _12263_/X _12269_/X VGND VGND VPWR VPWR _12747_/A sky130_fd_sc_hd__a21oi_4
XFILLER_107_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11221_ _11241_/A VGND VGND VPWR VPWR _11221_/X sky130_fd_sc_hd__buf_1
XFILLER_150_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11152_ _11518_/A VGND VGND VPWR VPWR _11152_/X sky130_fd_sc_hd__buf_1
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10103_ _14906_/Q _10097_/X _09969_/X _10098_/X VGND VGND VPWR VPWR _14906_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11083_ _11162_/A VGND VGND VPWR VPWR _11109_/A sky130_fd_sc_hd__buf_2
XFILLER_49_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14911_ _10083_/X _14911_/D VGND VGND VPWR VPWR _14911_/Q sky130_fd_sc_hd__dfxtp_1
X_10034_ _10403_/A VGND VGND VPWR VPWR _10034_/X sky130_fd_sc_hd__buf_1
XFILLER_102_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14842_ _10335_/X _14842_/D VGND VGND VPWR VPWR _14842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14773_ _10602_/X _14773_/D VGND VGND VPWR VPWR _14773_/Q sky130_fd_sc_hd__dfxtp_1
X_11985_ _11985_/A VGND VGND VPWR VPWR _12005_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10936_ _10936_/A VGND VGND VPWR VPWR _10936_/X sky130_fd_sc_hd__buf_1
XFILLER_32_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13724_ _15195_/Q _15163_/Q _14779_/Q _14811_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13724_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10867_ _10869_/A VGND VGND VPWR VPWR _10867_/X sky130_fd_sc_hd__clkbuf_1
X_13655_ _15138_/Q _15362_/Q _15330_/Q _15298_/Q _13740_/S0 _07541_/A VGND VGND VPWR
+ VPWR _13655_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12606_ _12065_/X _12602_/X _12829_/A VGND VGND VPWR VPWR _12606_/Y sky130_fd_sc_hd__o21ai_1
X_13586_ _13585_/X _14320_/D _15506_/Q VGND VGND VPWR VPWR _13586_/X sky130_fd_sc_hd__mux2_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10798_ _10798_/A VGND VGND VPWR VPWR _11541_/A sky130_fd_sc_hd__clkbuf_2
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15325_ _08381_/X _15325_/D VGND VGND VPWR VPWR _15325_/Q sky130_fd_sc_hd__dfxtp_1
X_12537_ _13162_/X _12493_/X _12525_/X _12528_/Y _12536_/X VGND VGND VPWR VPWR _12537_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_144_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15256_ _08706_/X _15256_/D VGND VGND VPWR VPWR _15256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12468_ _12435_/X _12440_/A _12443_/Y VGND VGND VPWR VPWR _12468_/X sky130_fd_sc_hd__o21a_1
X_11419_ _14566_/Q _11414_/X _11191_/X _11415_/X VGND VGND VPWR VPWR _14566_/D sky130_fd_sc_hd__a22o_1
X_14207_ _14635_/Q _14603_/Q _14571_/Q _15371_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14207_/X sky130_fd_sc_hd__mux4_1
X_15187_ _08983_/X _15187_/D VGND VGND VPWR VPWR _15187_/Q sky130_fd_sc_hd__dfxtp_1
X_12399_ _12371_/X _12381_/Y _12385_/X _12390_/X _12398_/X VGND VGND VPWR VPWR _12399_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_125_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14138_ _14514_/Q _14482_/Q _14450_/Q _14418_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14138_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14069_ _14841_/Q _14873_/Q _14905_/Q _14937_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14069_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_3_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR _14311_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08630_ _15277_/Q _08627_/X _08485_/X _08629_/X VGND VGND VPWR VPWR _15277_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08561_ _08574_/A VGND VGND VPWR VPWR _08572_/A sky130_fd_sc_hd__buf_1
XFILLER_70_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07512_ _07514_/A _07512_/B VGND VGND VPWR VPWR _15514_/D sky130_fd_sc_hd__nor2_1
XFILLER_35_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08492_ _09255_/A VGND VGND VPWR VPWR _08492_/X sky130_fd_sc_hd__buf_1
XFILLER_90_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07443_ _07443_/A VGND VGND VPWR VPWR _07446_/A sky130_fd_sc_hd__buf_1
XFILLER_90_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07374_ _07509_/B _07356_/X _12571_/A _07373_/X VGND VGND VPWR VPWR _07374_/X sky130_fd_sc_hd__o22a_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09113_ _15150_/Q _09106_/X _08873_/X _09107_/X VGND VGND VPWR VPWR _15150_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09044_ _09044_/A VGND VGND VPWR VPWR _09044_/X sky130_fd_sc_hd__buf_1
XFILLER_136_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09946_ _10026_/A VGND VGND VPWR VPWR _09974_/A sky130_fd_sc_hd__buf_2
X_09877_ _09877_/A VGND VGND VPWR VPWR _09877_/X sky130_fd_sc_hd__buf_1
X_08828_ _15225_/Q _08825_/X _08826_/X _08827_/X VGND VGND VPWR VPWR _15225_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08759_ _08761_/A VGND VGND VPWR VPWR _08759_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11770_ _14476_/Q _11764_/X _11533_/X _11766_/X VGND VGND VPWR VPWR _14476_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10721_ _10721_/A VGND VGND VPWR VPWR _10721_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13440_ _13696_/X _13701_/X _14386_/Q VGND VGND VPWR VPWR _13440_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10652_ _14758_/Q _10646_/X _10423_/X _10647_/X VGND VGND VPWR VPWR _14758_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13371_ _12610_/X _12577_/X _13418_/S VGND VGND VPWR VPWR _13371_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10583_ _10583_/A VGND VGND VPWR VPWR _10583_/X sky130_fd_sc_hd__buf_1
XFILLER_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12322_ _12456_/A VGND VGND VPWR VPWR _12878_/A sky130_fd_sc_hd__clkbuf_1
X_15110_ _09278_/X _15110_/D VGND VGND VPWR VPWR _15110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15041_ _09532_/X _15041_/D VGND VGND VPWR VPWR _15041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12253_ _12251_/X _12103_/A _12843_/A _12094_/X VGND VGND VPWR VPWR _12266_/B sky130_fd_sc_hd__o22a_1
XFILLER_108_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11204_ _11214_/A VGND VGND VPWR VPWR _11204_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12184_ _12274_/A _12183_/A _12752_/A _12183_/Y VGND VGND VPWR VPWR _12193_/A sky130_fd_sc_hd__o22a_1
XFILLER_69_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11135_ _11149_/A VGND VGND VPWR VPWR _11135_/X sky130_fd_sc_hd__buf_1
XFILLER_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11066_ _11078_/A VGND VGND VPWR VPWR _11082_/A sky130_fd_sc_hd__inv_2
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10017_ _14927_/Q _10011_/X _10016_/X _10013_/X VGND VGND VPWR VPWR _14927_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14825_ _10410_/X _14825_/D VGND VGND VPWR VPWR _14825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14756_ _10655_/X _14756_/D VGND VGND VPWR VPWR _14756_/Q sky130_fd_sc_hd__dfxtp_1
X_11968_ _14419_/Q _11966_/X _08016_/A _11967_/X VGND VGND VPWR VPWR _14419_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13707_ _14653_/Q _14621_/Q _14589_/Q _15389_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13707_/X sky130_fd_sc_hd__mux4_1
X_10919_ _14700_/Q _10914_/X _10788_/X _10916_/X VGND VGND VPWR VPWR _14700_/D sky130_fd_sc_hd__a22o_1
X_14687_ _10961_/X _14687_/D VGND VGND VPWR VPWR _14687_/Q sky130_fd_sc_hd__dfxtp_1
X_11899_ _14438_/Q _11895_/X _08084_/A _11896_/X VGND VGND VPWR VPWR _14438_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13638_ _13637_/X _14307_/D _15506_/Q VGND VGND VPWR VPWR _13638_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13569_ _13568_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13569_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15308_ _08489_/X _15308_/D VGND VGND VPWR VPWR _15308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15239_ _08761_/X _15239_/D VGND VGND VPWR VPWR _15239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09800_ _09802_/A VGND VGND VPWR VPWR _09800_/X sky130_fd_sc_hd__clkbuf_1
X_07992_ _08004_/A VGND VGND VPWR VPWR _07992_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09731_ _09731_/A VGND VGND VPWR VPWR _09731_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09662_ _10407_/A VGND VGND VPWR VPWR _09662_/X sky130_fd_sc_hd__buf_1
XFILLER_67_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08613_ _15281_/Q _08607_/X _08460_/X _08608_/X VGND VGND VPWR VPWR _15281_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09593_ _09625_/A VGND VGND VPWR VPWR _09593_/X sky130_fd_sc_hd__buf_1
XFILLER_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08544_ _10831_/A VGND VGND VPWR VPWR _09290_/A sky130_fd_sc_hd__buf_1
XFILLER_63_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08475_ _08489_/A VGND VGND VPWR VPWR _08475_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07426_ _07428_/A _13607_/X VGND VGND VPWR VPWR _15572_/D sky130_fd_sc_hd__and2_1
XFILLER_51_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07357_ _13648_/S VGND VGND VPWR VPWR _12574_/A sky130_fd_sc_hd__inv_2
XFILLER_108_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07288_ _07288_/A _07288_/B VGND VGND VPWR VPWR _15608_/D sky130_fd_sc_hd__nor2_1
XFILLER_108_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09027_ _15175_/Q _09025_/X _08905_/X _09026_/X VGND VGND VPWR VPWR _15175_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09929_ _09941_/A VGND VGND VPWR VPWR _09945_/A sky130_fd_sc_hd__inv_2
XFILLER_19_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12940_ _12708_/X _12712_/X _12914_/B _12939_/X VGND VGND VPWR VPWR _12941_/B sky130_fd_sc_hd__o22a_1
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12871_ _12670_/X _12869_/Y _12448_/X _12867_/Y _12870_/X VGND VGND VPWR VPWR _12871_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA_101 pc[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_112 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14610_ _11267_/X _14610_/D VGND VGND VPWR VPWR _14610_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_123 rdata[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 rdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11822_ _11828_/A VGND VGND VPWR VPWR _11822_/X sky130_fd_sc_hd__clkbuf_1
X_15590_ _15590_/CLK _15590_/D VGND VGND VPWR VPWR _15590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_145 rdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_167 wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11753_ _11753_/A VGND VGND VPWR VPWR _11753_/X sky130_fd_sc_hd__buf_1
XFILLER_26_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_178 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14541_ _11525_/X _14541_/D VGND VGND VPWR VPWR _14541_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_189 _12847_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10704_ _10719_/A VGND VGND VPWR VPWR _10704_/X sky130_fd_sc_hd__buf_1
XFILLER_42_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11684_ _14499_/Q _11578_/A _11570_/X _11581_/A VGND VGND VPWR VPWR _14499_/D sky130_fd_sc_hd__a22o_1
X_14472_ _11780_/X _14472_/D VGND VGND VPWR VPWR _14472_/Q sky130_fd_sc_hd__dfxtp_1
X_13423_ _12981_/X _12983_/Y _13425_/S VGND VGND VPWR VPWR _13423_/X sky130_fd_sc_hd__mux2_1
X_10635_ _14763_/Q _10627_/X _10403_/X _10629_/X VGND VGND VPWR VPWR _14763_/D sky130_fd_sc_hd__a22o_1
X_13354_ _12347_/X _12817_/B _15561_/Q VGND VGND VPWR VPWR _13354_/X sky130_fd_sc_hd__mux2_2
X_10566_ _10628_/A VGND VGND VPWR VPWR _10585_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12305_ _12307_/B VGND VGND VPWR VPWR _12324_/B sky130_fd_sc_hd__inv_2
X_13285_ _13284_/X _12323_/X _15565_/Q VGND VGND VPWR VPWR _13285_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10497_ _10506_/A VGND VGND VPWR VPWR _10497_/X sky130_fd_sc_hd__buf_1
X_15024_ _09624_/X _15024_/D VGND VGND VPWR VPWR _15024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12236_ _15568_/Q VGND VGND VPWR VPWR _12807_/A sky130_fd_sc_hd__inv_2
XFILLER_107_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12167_ _15541_/Q VGND VGND VPWR VPWR _12736_/A sky130_fd_sc_hd__buf_1
XFILLER_150_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11118_ _11125_/A VGND VGND VPWR VPWR _11118_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12098_ _12611_/A _12097_/A _12626_/A _12097_/Y VGND VGND VPWR VPWR _12580_/A sky130_fd_sc_hd__o22a_1
XFILLER_110_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11049_ _11049_/A VGND VGND VPWR VPWR _11054_/A sky130_fd_sc_hd__buf_1
XFILLER_110_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14808_ _10477_/X _14808_/D VGND VGND VPWR VPWR _14808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14739_ _10748_/X _14739_/D VGND VGND VPWR VPWR _14739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08260_ _08260_/A VGND VGND VPWR VPWR _08260_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07211_ _07247_/A VGND VGND VPWR VPWR _07246_/A sky130_fd_sc_hd__buf_1
X_08191_ _08191_/A VGND VGND VPWR VPWR _08264_/A sky130_fd_sc_hd__clkbuf_2
X_07142_ _13102_/X VGND VGND VPWR VPWR _07276_/B sky130_fd_sc_hd__inv_2
XFILLER_146_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07975_ _07975_/A VGND VGND VPWR VPWR _07986_/A sky130_fd_sc_hd__buf_1
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09714_ _09776_/A VGND VGND VPWR VPWR _09736_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09645_ _09678_/A VGND VGND VPWR VPWR _09645_/X sky130_fd_sc_hd__buf_1
XFILLER_71_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09576_ _09582_/A VGND VGND VPWR VPWR _09576_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _14307_/Q VGND VGND VPWR VPWR _10818_/A sky130_fd_sc_hd__buf_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _14318_/Q VGND VGND VPWR VPWR _10760_/A sky130_fd_sc_hd__buf_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ _07411_/A _13559_/X VGND VGND VPWR VPWR _15584_/D sky130_fd_sc_hd__and2_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08389_ _10702_/A VGND VGND VPWR VPWR _09184_/A sky130_fd_sc_hd__buf_1
XFILLER_7_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10420_ _10420_/A VGND VGND VPWR VPWR _10420_/X sky130_fd_sc_hd__buf_1
XFILLER_137_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10351_ _10358_/A VGND VGND VPWR VPWR _10351_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13070_ _12760_/Y _15572_/Q _13076_/S VGND VGND VPWR VPWR _13070_/X sky130_fd_sc_hd__mux2_1
X_10282_ _14855_/Q _10280_/X _10051_/X _10281_/X VGND VGND VPWR VPWR _14855_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12021_ _15585_/Q VGND VGND VPWR VPWR _12021_/X sky130_fd_sc_hd__buf_1
XFILLER_104_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13972_ _15234_/Q _14562_/Q _15010_/Q _15426_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13972_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12923_ _12805_/X _12235_/X _12806_/A _12807_/A VGND VGND VPWR VPWR _12933_/A sky130_fd_sc_hd__o22a_1
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15642_ _15648_/CLK _15642_/D VGND VGND VPWR VPWR _15642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12854_ _12854_/A VGND VGND VPWR VPWR _12854_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11805_ _11805_/A VGND VGND VPWR VPWR _11805_/X sky130_fd_sc_hd__clkbuf_1
X_15573_ _15667_/CLK _15573_/D VGND VGND VPWR VPWR _15573_/Q sky130_fd_sc_hd__dfxtp_1
X_12785_ _12785_/A _12785_/B _12847_/C VGND VGND VPWR VPWR _12785_/X sky130_fd_sc_hd__or3_1
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14524_ _11602_/X _14524_/D VGND VGND VPWR VPWR _14524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11736_ _14486_/Q _11733_/X _11489_/X _11735_/X VGND VGND VPWR VPWR _14486_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14455_ _11840_/X _14455_/D VGND VGND VPWR VPWR _14455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11667_ _11669_/A VGND VGND VPWR VPWR _11667_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _12635_/X _12634_/X _13418_/S VGND VGND VPWR VPWR _13406_/X sky130_fd_sc_hd__mux2_1
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10618_ _14768_/Q _10616_/X _10379_/X _10617_/X VGND VGND VPWR VPWR _14768_/D sky130_fd_sc_hd__a22o_1
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14386_ _14392_/CLK instruction[19] VGND VGND VPWR VPWR _14386_/Q sky130_fd_sc_hd__dfxtp_4
X_11598_ _11598_/A VGND VGND VPWR VPWR _11598_/X sky130_fd_sc_hd__clkbuf_1
X_13337_ _13383_/X _13381_/X _13415_/S VGND VGND VPWR VPWR _13337_/X sky130_fd_sc_hd__mux2_1
X_10549_ _10562_/A VGND VGND VPWR VPWR _10550_/A sky130_fd_sc_hd__buf_1
XFILLER_127_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13268_ _13269_/X _12878_/B _13393_/S VGND VGND VPWR VPWR _13268_/X sky130_fd_sc_hd__mux2_2
XFILLER_97_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15007_ _09712_/X _15007_/D VGND VGND VPWR VPWR _15007_/Q sky130_fd_sc_hd__dfxtp_1
X_12219_ _15563_/Q _12164_/X _12875_/A _12107_/A VGND VGND VPWR VPWR _12220_/A sky130_fd_sc_hd__o22a_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13199_ _13198_/X _12811_/X _15565_/Q VGND VGND VPWR VPWR _13199_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07760_ _13152_/X _07760_/B _07760_/C VGND VGND VPWR VPWR _07909_/B sky130_fd_sc_hd__or3_1
Xclkbuf_1_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_111_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07691_ _07653_/A _07686_/X _07695_/A _07690_/X VGND VGND VPWR VPWR _07779_/B sky130_fd_sc_hd__o211a_1
XFILLER_25_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09430_ _09439_/A VGND VGND VPWR VPWR _09435_/A sky130_fd_sc_hd__buf_1
XFILLER_18_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09361_ _09361_/A VGND VGND VPWR VPWR _09361_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08312_ _15340_/Q _08306_/X _08054_/X _08308_/X VGND VGND VPWR VPWR _15340_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09292_ _09307_/A VGND VGND VPWR VPWR _09305_/A sky130_fd_sc_hd__buf_1
XANTENNA_12 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08243_ _08307_/A VGND VGND VPWR VPWR _08262_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_34 data_address[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_45 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 instruction[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08174_ _08174_/A VGND VGND VPWR VPWR _08174_/X sky130_fd_sc_hd__buf_1
XANTENNA_78 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 pc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07125_ _13119_/X VGND VGND VPWR VPWR _07251_/B sky130_fd_sc_hd__inv_2
XFILLER_134_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07958_ _07958_/A VGND VGND VPWR VPWR _07958_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07889_ _07889_/A _07889_/B VGND VGND VPWR VPWR _07889_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09628_ _09628_/A VGND VGND VPWR VPWR _09628_/X sky130_fd_sc_hd__buf_1
XFILLER_16_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ _10324_/A VGND VGND VPWR VPWR _09559_/X sky130_fd_sc_hd__buf_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12570_ _12570_/A _12572_/B VGND VGND VPWR VPWR _12570_/X sky130_fd_sc_hd__or2_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ _11547_/A VGND VGND VPWR VPWR _11532_/A sky130_fd_sc_hd__buf_1
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240_ _14952_/Q _15048_/Q _15016_/Q _15080_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14240_/X sky130_fd_sc_hd__mux4_2
X_11452_ _11476_/A VGND VGND VPWR VPWR _11452_/X sky130_fd_sc_hd__buf_1
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10403_ _10403_/A VGND VGND VPWR VPWR _10403_/X sky130_fd_sc_hd__buf_1
X_14171_ _14167_/X _14168_/X _14169_/X _14170_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14171_/X sky130_fd_sc_hd__mux4_1
X_11383_ _11383_/A VGND VGND VPWR VPWR _11383_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13122_ _12492_/X _13025_/Y _13152_/S VGND VGND VPWR VPWR _13122_/X sky130_fd_sc_hd__mux2_2
X_10334_ _10334_/A VGND VGND VPWR VPWR _10343_/A sky130_fd_sc_hd__clkbuf_2
X_13053_ wdata[26] rdata[26] _13057_/S VGND VGND VPWR VPWR _14330_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10265_ _14859_/Q _10257_/X _10034_/X _10259_/X VGND VGND VPWR VPWR _14859_/D sky130_fd_sc_hd__a22o_1
XFILLER_140_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12004_ _12010_/A VGND VGND VPWR VPWR _12004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10196_ _10217_/A VGND VGND VPWR VPWR _10196_/X sky130_fd_sc_hd__buf_1
XFILLER_66_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13955_ _15108_/Q _15332_/Q _15300_/Q _15268_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13955_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12906_ _12946_/C _12906_/B VGND VGND VPWR VPWR _12909_/C sky130_fd_sc_hd__or2_1
XFILLER_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13886_ _13882_/X _13883_/X _13884_/X _13885_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13886_/X sky130_fd_sc_hd__mux4_2
XFILLER_46_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15625_ _15654_/CLK _15625_/D VGND VGND VPWR VPWR pc[20] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12837_ _12837_/A VGND VGND VPWR VPWR _12838_/A sky130_fd_sc_hd__buf_1
XFILLER_15_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15556_ _15589_/CLK _15556_/D VGND VGND VPWR VPWR _15556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12768_ _12749_/A _12749_/B _12512_/X _12750_/B VGND VGND VPWR VPWR _12768_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14507_ _11658_/X _14507_/D VGND VGND VPWR VPWR _14507_/Q sky130_fd_sc_hd__dfxtp_1
X_11719_ _11721_/A VGND VGND VPWR VPWR _11719_/X sky130_fd_sc_hd__clkbuf_1
X_15487_ _15667_/CLK _15487_/D VGND VGND VPWR VPWR wdata[13] sky130_fd_sc_hd__dfxtp_4
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12699_ _12699_/A _12699_/B VGND VGND VPWR VPWR _12783_/A sky130_fd_sc_hd__or2_1
XFILLER_30_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14438_ _11898_/X _14438_/D VGND VGND VPWR VPWR _14438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14369_ _14392_/CLK pc[30] VGND VGND VPWR VPWR _14369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08930_ _08941_/A VGND VGND VPWR VPWR _08944_/A sky130_fd_sc_hd__inv_2
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08861_ _09232_/A VGND VGND VPWR VPWR _08861_/X sky130_fd_sc_hd__buf_1
XFILLER_69_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07812_ _07805_/A _07805_/B _07796_/X _07805_/Y VGND VGND VPWR VPWR _15453_/D sky130_fd_sc_hd__o211a_1
X_08792_ _08804_/A VGND VGND VPWR VPWR _08792_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07743_ _13146_/X VGND VGND VPWR VPWR _07743_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07674_ _13128_/X VGND VGND VPWR VPWR _07674_/X sky130_fd_sc_hd__buf_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09413_ _09413_/A VGND VGND VPWR VPWR _09413_/X sky130_fd_sc_hd__buf_1
XFILLER_41_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09344_ _09374_/A VGND VGND VPWR VPWR _09365_/A sky130_fd_sc_hd__buf_2
X_09275_ _09275_/A VGND VGND VPWR VPWR _09275_/X sky130_fd_sc_hd__buf_1
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08226_ _08239_/A VGND VGND VPWR VPWR _08227_/A sky130_fd_sc_hd__buf_1
XFILLER_147_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08157_ _08159_/A VGND VGND VPWR VPWR _08157_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07108_ _07586_/A VGND VGND VPWR VPWR _07795_/A sky130_fd_sc_hd__buf_1
X_08088_ _08118_/A VGND VGND VPWR VPWR _08097_/A sky130_fd_sc_hd__buf_1
XFILLER_106_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10050_ _10050_/A VGND VGND VPWR VPWR _10050_/X sky130_fd_sc_hd__buf_1
XFILLER_87_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13740_ _14970_/Q _15066_/Q _15034_/Q _15098_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13740_/X sky130_fd_sc_hd__mux4_2
X_10952_ _10962_/A VGND VGND VPWR VPWR _10965_/A sky130_fd_sc_hd__inv_2
XFILLER_44_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13671_ _13667_/X _13668_/X _13669_/X _13670_/X _07533_/A _14402_/Q VGND VGND VPWR
+ VPWR _13671_/X sky130_fd_sc_hd__mux4_1
X_10883_ _10913_/A VGND VGND VPWR VPWR _10904_/A sky130_fd_sc_hd__buf_1
XFILLER_71_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15410_ _08019_/X _15410_/D VGND VGND VPWR VPWR _15410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12622_ _12946_/C VGND VGND VPWR VPWR _12622_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15341_ _08304_/X _15341_/D VGND VGND VPWR VPWR _15341_/Q sky130_fd_sc_hd__dfxtp_1
X_12553_ _12553_/A VGND VGND VPWR VPWR _12553_/X sky130_fd_sc_hd__buf_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11504_ _14547_/Q _11501_/X _11502_/X _11503_/X VGND VGND VPWR VPWR _14547_/D sky130_fd_sc_hd__a22o_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15272_ _08642_/X _15272_/D VGND VGND VPWR VPWR _15272_/Q sky130_fd_sc_hd__dfxtp_1
X_12484_ _12819_/A VGND VGND VPWR VPWR _12770_/A sky130_fd_sc_hd__clkbuf_1
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14223_ _14665_/Q _15241_/Q _14729_/Q _14697_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14223_/X sky130_fd_sc_hd__mux4_2
X_11435_ _14562_/Q _11430_/X _11431_/X _11434_/X VGND VGND VPWR VPWR _14562_/D sky130_fd_sc_hd__a22o_1
XFILLER_153_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14154_ _15184_/Q _15152_/Q _14768_/Q _14800_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14154_/X sky130_fd_sc_hd__mux4_1
X_11366_ _11385_/A VGND VGND VPWR VPWR _11366_/X sky130_fd_sc_hd__buf_1
XFILLER_125_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13105_ _15651_/Q data_address[16] _15667_/Q VGND VGND VPWR VPWR _13105_/X sky130_fd_sc_hd__mux2_1
X_10317_ _10341_/A VGND VGND VPWR VPWR _10317_/X sky130_fd_sc_hd__buf_1
X_11297_ _11299_/A VGND VGND VPWR VPWR _11297_/X sky130_fd_sc_hd__clkbuf_1
X_14085_ _15127_/Q _15351_/Q _15319_/Q _15287_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14085_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10248_ _10248_/A VGND VGND VPWR VPWR _10248_/X sky130_fd_sc_hd__buf_1
X_13036_ wdata[9] rdata[9] _13057_/S VGND VGND VPWR VPWR _14313_/D sky130_fd_sc_hd__mux2_2
XFILLER_94_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10179_ _14883_/Q _10071_/A _10065_/X _10074_/A VGND VGND VPWR VPWR _14883_/D sky130_fd_sc_hd__a22o_1
XFILLER_121_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14987_ _09783_/X _14987_/D VGND VGND VPWR VPWR _14987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13938_ _14502_/Q _14470_/Q _14438_/Q _14406_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13938_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13869_ _14829_/Q _14861_/Q _14893_/Q _14925_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13869_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15608_ _15648_/CLK _15608_/D VGND VGND VPWR VPWR pc[3] sky130_fd_sc_hd__dfxtp_1
X_07390_ _07386_/Y _07363_/A _07510_/B _07319_/A _07389_/X VGND VGND VPWR VPWR _07392_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_50_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15539_ _15576_/CLK _15539_/D VGND VGND VPWR VPWR _15539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09060_ _09064_/A VGND VGND VPWR VPWR _09060_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08011_ _08011_/A VGND VGND VPWR VPWR _08011_/X sky130_fd_sc_hd__buf_1
XFILLER_129_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09962_ _10332_/A VGND VGND VPWR VPWR _09962_/X sky130_fd_sc_hd__buf_1
X_08913_ _09284_/A VGND VGND VPWR VPWR _08913_/X sky130_fd_sc_hd__buf_1
XFILLER_69_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09893_ _09897_/A VGND VGND VPWR VPWR _09893_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08844_ _09216_/A VGND VGND VPWR VPWR _08844_/X sky130_fd_sc_hd__buf_1
XFILLER_111_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08775_ _08788_/A VGND VGND VPWR VPWR _08775_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07726_ _07723_/X _07725_/X _13142_/X _07725_/A VGND VGND VPWR VPWR _07873_/A sky130_fd_sc_hd__a2bb2o_1
X_07657_ _07786_/A VGND VGND VPWR VPWR _07658_/A sky130_fd_sc_hd__buf_1
XFILLER_13_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07588_ _07596_/A VGND VGND VPWR VPWR _07591_/A sky130_fd_sc_hd__buf_1
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09327_ _09336_/A VGND VGND VPWR VPWR _09327_/X sky130_fd_sc_hd__buf_1
XFILLER_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09258_ _09266_/A VGND VGND VPWR VPWR _09258_/X sky130_fd_sc_hd__clkbuf_1
X_08209_ _08209_/A VGND VGND VPWR VPWR _08209_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09189_ _15131_/Q _09183_/X _09188_/X _09185_/X VGND VGND VPWR VPWR _15131_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11220_ _11283_/A VGND VGND VPWR VPWR _11241_/A sky130_fd_sc_hd__buf_2
XFILLER_153_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11151_ _11151_/A VGND VGND VPWR VPWR _11151_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10102_ _10102_/A VGND VGND VPWR VPWR _10102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11082_ _11082_/A VGND VGND VPWR VPWR _11162_/A sky130_fd_sc_hd__buf_2
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10033_ _10041_/A VGND VGND VPWR VPWR _10033_/X sky130_fd_sc_hd__clkbuf_1
X_14910_ _10091_/X _14910_/D VGND VGND VPWR VPWR _14910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14841_ _10338_/X _14841_/D VGND VGND VPWR VPWR _14841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14772_ _10604_/X _14772_/D VGND VGND VPWR VPWR _14772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11984_ _11992_/A VGND VGND VPWR VPWR _11984_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13723_ _14683_/Q _15259_/Q _14747_/Q _14715_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13723_/X sky130_fd_sc_hd__mux4_2
X_10935_ _10941_/A VGND VGND VPWR VPWR _10935_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13654_ _15202_/Q _15170_/Q _14786_/Q _14818_/Q _13740_/S0 _07541_/A VGND VGND VPWR
+ VPWR _13654_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10866_ _14716_/Q _10864_/X _10703_/X _10865_/X VGND VGND VPWR VPWR _14716_/D sky130_fd_sc_hd__a22o_1
XFILLER_16_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12605_ _12605_/A VGND VGND VPWR VPWR _12829_/A sky130_fd_sc_hd__buf_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _13584_/X _07310_/Y _13649_/S VGND VGND VPWR VPWR _13585_/X sky130_fd_sc_hd__mux2_1
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10797_ _10812_/A VGND VGND VPWR VPWR _10797_/X sky130_fd_sc_hd__buf_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15324_ _08386_/X _15324_/D VGND VGND VPWR VPWR _15324_/Q sky130_fd_sc_hd__dfxtp_1
X_12536_ _12530_/Y _12534_/A _12530_/A _12534_/Y _12535_/X VGND VGND VPWR VPWR _12536_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15255_ _08708_/X _15255_/D VGND VGND VPWR VPWR _15255_/Q sky130_fd_sc_hd__dfxtp_1
X_12467_ _12509_/A _12509_/B _12466_/Y VGND VGND VPWR VPWR _12467_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_8_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14206_ _14202_/X _14203_/X _14204_/X _14205_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14206_/X sky130_fd_sc_hd__mux4_2
XFILLER_144_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11418_ _11422_/A VGND VGND VPWR VPWR _11418_/X sky130_fd_sc_hd__clkbuf_1
X_15186_ _08987_/X _15186_/D VGND VGND VPWR VPWR _15186_/Q sky130_fd_sc_hd__dfxtp_1
X_12398_ _12432_/A _12397_/B _12578_/A _12410_/B VGND VGND VPWR VPWR _12398_/X sky130_fd_sc_hd__a211o_1
XFILLER_99_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14137_ _14642_/Q _14610_/Q _14578_/Q _15378_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14137_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11349_ _11353_/A VGND VGND VPWR VPWR _11349_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14068_ _14521_/Q _14489_/Q _14457_/Q _14425_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14068_/X sky130_fd_sc_hd__mux4_2
XFILLER_95_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13019_ _14363_/Q VGND VGND VPWR VPWR _13019_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08560_ _15296_/Q _08552_/X _08361_/X _08555_/X VGND VGND VPWR VPWR _15296_/D sky130_fd_sc_hd__a22o_1
X_07511_ _07511_/A VGND VGND VPWR VPWR _07514_/A sky130_fd_sc_hd__buf_1
X_08491_ _10787_/A VGND VGND VPWR VPWR _09255_/A sky130_fd_sc_hd__buf_1
XFILLER_35_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07442_ _07442_/A _13651_/X VGND VGND VPWR VPWR _15561_/D sky130_fd_sc_hd__and2_1
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07373_ _07373_/A VGND VGND VPWR VPWR _07373_/X sky130_fd_sc_hd__buf_1
XFILLER_148_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09112_ _09114_/A VGND VGND VPWR VPWR _09112_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09043_ _09055_/A VGND VGND VPWR VPWR _09044_/A sky130_fd_sc_hd__buf_1
XFILLER_135_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09945_ _09945_/A VGND VGND VPWR VPWR _10026_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09876_ _09876_/A VGND VGND VPWR VPWR _09876_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08827_ _08827_/A VGND VGND VPWR VPWR _08827_/X sky130_fd_sc_hd__buf_1
XFILLER_85_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08758_ _15241_/Q _08753_/X _08511_/X _08754_/X VGND VGND VPWR VPWR _15241_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07709_ _13140_/X VGND VGND VPWR VPWR _07709_/X sky130_fd_sc_hd__buf_1
XFILLER_72_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08689_ _15262_/Q _08679_/X _08377_/X _08682_/X VGND VGND VPWR VPWR _15262_/D sky130_fd_sc_hd__a22o_1
XFILLER_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10720_ _14745_/Q _10716_/X _10718_/X _10719_/X VGND VGND VPWR VPWR _14745_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10651_ _10655_/A VGND VGND VPWR VPWR _10651_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13370_ _12590_/X _12329_/X _13418_/S VGND VGND VPWR VPWR _13370_/X sky130_fd_sc_hd__mux2_1
X_10582_ _14778_/Q _10575_/X _10336_/X _10576_/X VGND VGND VPWR VPWR _14778_/D sky130_fd_sc_hd__a22o_1
X_12321_ _12343_/A VGND VGND VPWR VPWR _12456_/A sky130_fd_sc_hd__buf_1
XFILLER_108_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15040_ _09537_/X _15040_/D VGND VGND VPWR VPWR _15040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12252_ _15566_/Q VGND VGND VPWR VPWR _12843_/A sky130_fd_sc_hd__inv_2
XFILLER_123_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11203_ _11203_/A VGND VGND VPWR VPWR _11214_/A sky130_fd_sc_hd__buf_1
X_12183_ _12183_/A VGND VGND VPWR VPWR _12183_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11134_ _11502_/A VGND VGND VPWR VPWR _11134_/X sky130_fd_sc_hd__buf_1
XFILLER_122_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11065_ _11431_/A VGND VGND VPWR VPWR _11065_/X sky130_fd_sc_hd__buf_1
XFILLER_89_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10016_ _10383_/A VGND VGND VPWR VPWR _10016_/X sky130_fd_sc_hd__buf_1
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14824_ _10414_/X _14824_/D VGND VGND VPWR VPWR _14824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14755_ _10658_/X _14755_/D VGND VGND VPWR VPWR _14755_/Q sky130_fd_sc_hd__dfxtp_1
X_11967_ _11977_/A VGND VGND VPWR VPWR _11967_/X sky130_fd_sc_hd__buf_1
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13706_ _13702_/X _13703_/X _13704_/X _13705_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13706_/X sky130_fd_sc_hd__mux4_2
X_10918_ _10920_/A VGND VGND VPWR VPWR _10918_/X sky130_fd_sc_hd__clkbuf_1
X_14686_ _10971_/X _14686_/D VGND VGND VPWR VPWR _14686_/Q sky130_fd_sc_hd__dfxtp_1
X_11898_ _11898_/A VGND VGND VPWR VPWR _11898_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13637_ _13636_/X _07369_/Y _13641_/S VGND VGND VPWR VPWR _13637_/X sky130_fd_sc_hd__mux2_1
X_10849_ _10862_/A VGND VGND VPWR VPWR _10860_/A sky130_fd_sc_hd__buf_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13568_ _14086_/X _14091_/X _13648_/S VGND VGND VPWR VPWR _13568_/X sky130_fd_sc_hd__mux2_1
X_15307_ _08496_/X _15307_/D VGND VGND VPWR VPWR _15307_/Q sky130_fd_sc_hd__dfxtp_1
X_12519_ _12519_/A _12519_/B VGND VGND VPWR VPWR _12520_/B sky130_fd_sc_hd__or2_1
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13499_ _13498_/X _13067_/X _14336_/Q VGND VGND VPWR VPWR _13499_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15238_ _08766_/X _15238_/D VGND VGND VPWR VPWR _15238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15169_ _09047_/X _15169_/D VGND VGND VPWR VPWR _15169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07991_ _08023_/A VGND VGND VPWR VPWR _08004_/A sky130_fd_sc_hd__buf_1
XFILLER_68_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09730_ _15003_/Q _09726_/X _09569_/X _09727_/X VGND VGND VPWR VPWR _15003_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09661_ _10798_/A VGND VGND VPWR VPWR _10407_/A sky130_fd_sc_hd__buf_1
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08612_ _08612_/A VGND VGND VPWR VPWR _08612_/X sky130_fd_sc_hd__clkbuf_1
X_09592_ _09640_/A VGND VGND VPWR VPWR _09625_/A sky130_fd_sc_hd__buf_2
XFILLER_36_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08543_ _14304_/Q VGND VGND VPWR VPWR _10831_/A sky130_fd_sc_hd__buf_1
XFILLER_70_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08474_ _08474_/A VGND VGND VPWR VPWR _08489_/A sky130_fd_sc_hd__buf_2
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07425_ _07429_/A VGND VGND VPWR VPWR _07428_/A sky130_fd_sc_hd__clkbuf_1
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07356_ _07356_/A VGND VGND VPWR VPWR _07356_/X sky130_fd_sc_hd__buf_1
X_07287_ _07288_/A _07287_/B VGND VGND VPWR VPWR _15609_/D sky130_fd_sc_hd__nor2_1
X_09026_ _09026_/A VGND VGND VPWR VPWR _09026_/X sky130_fd_sc_hd__buf_1
XFILLER_105_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09928_ _10297_/A VGND VGND VPWR VPWR _09928_/X sky130_fd_sc_hd__buf_1
XFILLER_19_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09859_ _14966_/Q _09856_/X _09595_/X _09858_/X VGND VGND VPWR VPWR _14966_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12870_ _12213_/Y _12211_/X _12336_/A _13327_/X _12741_/X VGND VGND VPWR VPWR _12870_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_65_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_102 pc[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_113 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11821_ _11839_/A VGND VGND VPWR VPWR _11828_/A sky130_fd_sc_hd__buf_1
XFILLER_61_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_124 rdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_135 rdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_146 rdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_157 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14540_ _11532_/X _14540_/D VGND VGND VPWR VPWR _14540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11752_ _11752_/A VGND VGND VPWR VPWR _11752_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_168 wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_179 wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10703_ _11463_/A VGND VGND VPWR VPWR _10703_/X sky130_fd_sc_hd__buf_1
X_14471_ _11782_/X _14471_/D VGND VGND VPWR VPWR _14471_/Q sky130_fd_sc_hd__dfxtp_1
X_11683_ _11685_/A VGND VGND VPWR VPWR _11683_/X sky130_fd_sc_hd__clkbuf_1
X_13422_ _12029_/Y _12052_/X _13425_/S VGND VGND VPWR VPWR _13422_/X sky130_fd_sc_hd__mux2_1
X_10634_ _10636_/A VGND VGND VPWR VPWR _10634_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13353_ _13416_/X _13414_/X _13415_/S VGND VGND VPWR VPWR _13353_/X sky130_fd_sc_hd__mux2_1
X_10565_ _10565_/A VGND VGND VPWR VPWR _10628_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_127_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12304_ _12329_/A _12303_/B _12357_/A VGND VGND VPWR VPWR _12431_/A sky130_fd_sc_hd__a21o_1
XFILLER_127_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13284_ _13408_/X _13401_/X _13393_/S VGND VGND VPWR VPWR _13284_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10496_ _10505_/A VGND VGND VPWR VPWR _10496_/X sky130_fd_sc_hd__buf_1
XFILLER_6_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15023_ _09630_/X _15023_/D VGND VGND VPWR VPWR _15023_/Q sky130_fd_sc_hd__dfxtp_1
X_12235_ _15568_/Q VGND VGND VPWR VPWR _12235_/X sky130_fd_sc_hd__buf_1
XFILLER_142_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12166_ _15573_/Q _12164_/X _12737_/B _12130_/X VGND VGND VPWR VPWR _12168_/A sky130_fd_sc_hd__o22a_1
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11117_ _14647_/Q _11107_/X _11116_/X _11109_/X VGND VGND VPWR VPWR _14647_/D sky130_fd_sc_hd__a22o_1
X_12097_ _12097_/A VGND VGND VPWR VPWR _12097_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11048_ _14663_/Q _11046_/X _10814_/X _11047_/X VGND VGND VPWR VPWR _14663_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14807_ _10479_/X _14807_/D VGND VGND VPWR VPWR _14807_/Q sky130_fd_sc_hd__dfxtp_1
X_12999_ _14343_/Q VGND VGND VPWR VPWR _12999_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14738_ _10754_/X _14738_/D VGND VGND VPWR VPWR _14738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14669_ _11023_/X _14669_/D VGND VGND VPWR VPWR _14669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07210_ _13108_/X _07208_/Y _07209_/X _07169_/B VGND VGND VPWR VPWR _15654_/D sky130_fd_sc_hd__o211a_1
X_08190_ _15371_/Q _08183_/X _08059_/X _08185_/X VGND VGND VPWR VPWR _15371_/D sky130_fd_sc_hd__a22o_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07141_ _13103_/X VGND VGND VPWR VPWR _07273_/B sky130_fd_sc_hd__inv_2
XFILLER_146_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_opt_9_clk _14328_/CLK VGND VGND VPWR VPWR _14324_/CLK sky130_fd_sc_hd__clkbuf_16
X_07974_ _15419_/Q _07966_/X _07973_/X _07969_/X VGND VGND VPWR VPWR _15419_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09713_ _09713_/A VGND VGND VPWR VPWR _09776_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09644_ _09644_/A VGND VGND VPWR VPWR _09678_/A sky130_fd_sc_hd__buf_1
XFILLER_83_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09575_ _15034_/Q _09562_/X _09574_/X _09565_/X VGND VGND VPWR VPWR _15034_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08526_ _08526_/A VGND VGND VPWR VPWR _08526_/X sky130_fd_sc_hd__clkbuf_1
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08457_ _08469_/A VGND VGND VPWR VPWR _08457_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07408_ _07416_/A VGND VGND VPWR VPWR _07411_/A sky130_fd_sc_hd__buf_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08388_ _14329_/Q VGND VGND VPWR VPWR _10702_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07339_ _07354_/A VGND VGND VPWR VPWR _07339_/X sky130_fd_sc_hd__buf_1
X_10350_ _14839_/Q _10339_/X _10349_/X _10341_/X VGND VGND VPWR VPWR _14839_/D sky130_fd_sc_hd__a22o_1
XFILLER_137_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09009_ _15181_/Q _09006_/X _08878_/X _09008_/X VGND VGND VPWR VPWR _15181_/D sky130_fd_sc_hd__a22o_1
X_10281_ _10281_/A VGND VGND VPWR VPWR _10281_/X sky130_fd_sc_hd__buf_1
XFILLER_151_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12020_ _15553_/Q VGND VGND VPWR VPWR _12020_/X sky130_fd_sc_hd__buf_1
XFILLER_105_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13971_ _13967_/X _13968_/X _13969_/X _13970_/X _07533_/A _14402_/Q VGND VGND VPWR
+ VPWR _13971_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12922_ _12828_/X _12243_/X _12820_/A _12825_/A VGND VGND VPWR VPWR _12924_/C sky130_fd_sc_hd__o22a_1
XFILLER_19_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15641_ _15648_/CLK _15641_/D VGND VGND VPWR VPWR _15641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12853_ _12852_/X _12838_/X _12789_/X _13318_/X _12826_/X VGND VGND VPWR VPWR _12853_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11804_ _14466_/Q _11800_/X _07929_/A _11803_/X VGND VGND VPWR VPWR _14466_/D sky130_fd_sc_hd__a22o_1
X_15572_ _15576_/CLK _15572_/D VGND VGND VPWR VPWR _15572_/Q sky130_fd_sc_hd__dfxtp_1
X_12784_ _12784_/A VGND VGND VPWR VPWR _12847_/C sky130_fd_sc_hd__clkbuf_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14523_ _11606_/X _14523_/D VGND VGND VPWR VPWR _14523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11735_ _11753_/A VGND VGND VPWR VPWR _11735_/X sky130_fd_sc_hd__buf_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14454_ _11842_/X _14454_/D VGND VGND VPWR VPWR _14454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11666_ _14506_/Q _11664_/X _11541_/X _11665_/X VGND VGND VPWR VPWR _14506_/D sky130_fd_sc_hd__a22o_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _13407_/X _13406_/X _13415_/S VGND VGND VPWR VPWR _13405_/X sky130_fd_sc_hd__mux2_1
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10617_ _10617_/A VGND VGND VPWR VPWR _10617_/X sky130_fd_sc_hd__buf_1
Xclkbuf_opt_10_clk _14328_/CLK VGND VGND VPWR VPWR _14379_/CLK sky130_fd_sc_hd__clkbuf_16
X_14385_ _14385_/CLK instruction[14] VGND VGND VPWR VPWR _14385_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11597_ _14526_/Q _11591_/X _11455_/X _11594_/X VGND VGND VPWR VPWR _14526_/D sky130_fd_sc_hd__a22o_1
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13336_ _13380_/X _13378_/X _13415_/S VGND VGND VPWR VPWR _13336_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10548_ _10548_/A _10548_/B VGND VGND VPWR VPWR _10562_/A sky130_fd_sc_hd__or2_2
XFILLER_115_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13267_ _13266_/X _12400_/X _15565_/Q VGND VGND VPWR VPWR _13267_/X sky130_fd_sc_hd__mux2_1
X_10479_ _10479_/A VGND VGND VPWR VPWR _10479_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15006_ _09720_/X _15006_/D VGND VGND VPWR VPWR _15006_/Q sky130_fd_sc_hd__dfxtp_1
X_12218_ _15563_/Q VGND VGND VPWR VPWR _12875_/A sky130_fd_sc_hd__inv_2
X_13198_ _13200_/X _13239_/X _13393_/S VGND VGND VPWR VPWR _13198_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12149_ _12146_/X _12164_/A _12694_/A _12148_/X VGND VGND VPWR VPWR _12150_/A sky130_fd_sc_hd__o22a_1
XFILLER_96_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07690_ _07682_/X _07688_/X _07689_/X _13129_/X VGND VGND VPWR VPWR _07690_/X sky130_fd_sc_hd__o22a_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09360_ _15090_/Q _09356_/X _09228_/X _09357_/X VGND VGND VPWR VPWR _15090_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08311_ _08315_/A VGND VGND VPWR VPWR _08311_/X sky130_fd_sc_hd__clkbuf_1
X_09291_ _15107_/Q _09152_/A _09290_/X _09156_/A VGND VGND VPWR VPWR _15107_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08242_ _08242_/A VGND VGND VPWR VPWR _08307_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_24 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_35 data_address[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08173_ _08173_/A VGND VGND VPWR VPWR _08173_/X sky130_fd_sc_hd__buf_1
XANTENNA_68 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 pc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07124_ _07820_/A _13059_/X _13152_/S VGND VGND VPWR VPWR _15667_/D sky130_fd_sc_hd__and3_1
XFILLER_118_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07957_ _14331_/Q VGND VGND VPWR VPWR _07958_/A sky130_fd_sc_hd__buf_1
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07888_ _07884_/A _07884_/B _07882_/X _07885_/A VGND VGND VPWR VPWR _15435_/D sky130_fd_sc_hd__o211a_1
XFILLER_16_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09627_ _10379_/A VGND VGND VPWR VPWR _09627_/X sky130_fd_sc_hd__buf_1
XFILLER_71_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09558_ _10697_/A VGND VGND VPWR VPWR _10324_/A sky130_fd_sc_hd__buf_1
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08509_ _14310_/Q VGND VGND VPWR VPWR _10803_/A sky130_fd_sc_hd__buf_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09489_ _15053_/Q _09486_/X _09250_/X _09488_/X VGND VGND VPWR VPWR _15053_/D sky130_fd_sc_hd__a22o_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _11520_/A VGND VGND VPWR VPWR _11547_/A sky130_fd_sc_hd__buf_1
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11451_ _11529_/A VGND VGND VPWR VPWR _11476_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10402_ _10410_/A VGND VGND VPWR VPWR _10402_/X sky130_fd_sc_hd__clkbuf_1
X_14170_ _14959_/Q _15055_/Q _15023_/Q _15087_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14170_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11382_ _14577_/Q _11374_/X _11144_/X _11375_/X VGND VGND VPWR VPWR _14577_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13121_ _15560_/Q _14370_/Q _13152_/S VGND VGND VPWR VPWR _13121_/X sky130_fd_sc_hd__mux2_1
X_10333_ _14843_/Q _10327_/X _10332_/X _10329_/X VGND VGND VPWR VPWR _14843_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13052_ wdata[25] rdata[25] _13057_/S VGND VGND VPWR VPWR _14329_/D sky130_fd_sc_hd__mux2_1
X_10264_ _10266_/A VGND VGND VPWR VPWR _10264_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12003_ _12012_/A VGND VGND VPWR VPWR _12010_/A sky130_fd_sc_hd__buf_1
XFILLER_133_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10195_ _10256_/A VGND VGND VPWR VPWR _10217_/A sky130_fd_sc_hd__buf_2
XFILLER_120_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13954_ _15172_/Q _15140_/Q _14756_/Q _14788_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13954_/X sky130_fd_sc_hd__mux4_1
X_12905_ _12905_/A _12905_/B _12905_/C VGND VGND VPWR VPWR _12959_/C sky130_fd_sc_hd__or3_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13885_ _15115_/Q _15339_/Q _15307_/Q _15275_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13885_/X sky130_fd_sc_hd__mux4_2
X_15624_ _15654_/CLK _15624_/D VGND VGND VPWR VPWR pc[19] sky130_fd_sc_hd__dfxtp_1
X_12836_ _12836_/A VGND VGND VPWR VPWR _12847_/A sky130_fd_sc_hd__buf_4
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15555_ _15589_/CLK _15555_/D VGND VGND VPWR VPWR _15555_/Q sky130_fd_sc_hd__dfxtp_1
X_12767_ _12765_/X _12187_/X _12713_/X _12766_/X VGND VGND VPWR VPWR _12767_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_70_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14506_ _11663_/X _14506_/D VGND VGND VPWR VPWR _14506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11718_ _14491_/Q _11713_/X _11467_/X _11714_/X VGND VGND VPWR VPWR _14491_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15486_ _15667_/CLK _15486_/D VGND VGND VPWR VPWR wdata[12] sky130_fd_sc_hd__dfxtp_1
X_12698_ _12826_/A VGND VGND VPWR VPWR _12698_/X sky130_fd_sc_hd__buf_1
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14437_ _11901_/X _14437_/D VGND VGND VPWR VPWR _14437_/Q sky130_fd_sc_hd__dfxtp_1
X_11649_ _11649_/A VGND VGND VPWR VPWR _11658_/A sky130_fd_sc_hd__buf_1
XFILLER_128_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14368_ _15666_/CLK pc[29] VGND VGND VPWR VPWR _14368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13319_ _13320_/X _12425_/B _13393_/S VGND VGND VPWR VPWR _13319_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14299_ _15469_/CLK _15466_/Q VGND VGND VPWR VPWR _14299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08860_ _08868_/A VGND VGND VPWR VPWR _08860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07811_ _07808_/A _07807_/Y _07808_/Y _07807_/A _07810_/X VGND VGND VPWR VPWR _15454_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08791_ _08807_/A VGND VGND VPWR VPWR _08804_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07742_ _15599_/Q VGND VGND VPWR VPWR _07742_/Y sky130_fd_sc_hd__inv_2
X_07673_ _07655_/A _13125_/X _07655_/A _13125_/X VGND VGND VPWR VPWR _07808_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09412_ _09426_/A VGND VGND VPWR VPWR _09413_/A sky130_fd_sc_hd__buf_1
XFILLER_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09343_ _09351_/A VGND VGND VPWR VPWR _09343_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09274_ _09274_/A VGND VGND VPWR VPWR _09274_/X sky130_fd_sc_hd__buf_1
XFILLER_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08225_ _09150_/A _11686_/A VGND VGND VPWR VPWR _08239_/A sky130_fd_sc_hd__or2_2
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08156_ _15382_/Q _08153_/X _08000_/X _08155_/X VGND VGND VPWR VPWR _15382_/D sky130_fd_sc_hd__a22o_1
X_07107_ _15667_/Q VGND VGND VPWR VPWR _07586_/A sky130_fd_sc_hd__inv_2
XFILLER_134_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08087_ _08161_/A VGND VGND VPWR VPWR _08118_/A sky130_fd_sc_hd__buf_2
XFILLER_103_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08989_ _08989_/A VGND VGND VPWR VPWR _08989_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10951_ _10951_/A VGND VGND VPWR VPWR _10951_/X sky130_fd_sc_hd__buf_1
XFILLER_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13670_ _14977_/Q _15073_/Q _15041_/Q _15105_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13670_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10882_ _10890_/A VGND VGND VPWR VPWR _10882_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12621_ _12615_/X _12101_/X _12610_/X _12618_/X VGND VGND VPWR VPWR _12946_/C sky130_fd_sc_hd__o22a_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15340_ _08311_/X _15340_/D VGND VGND VPWR VPWR _15340_/Q sky130_fd_sc_hd__dfxtp_1
X_12552_ _12545_/A _12550_/Y _12545_/C _12551_/Y _12541_/B VGND VGND VPWR VPWR _12553_/A
+ sky130_fd_sc_hd__o221a_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _11515_/A VGND VGND VPWR VPWR _11503_/X sky130_fd_sc_hd__buf_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15271_ _08646_/X _15271_/D VGND VGND VPWR VPWR _15271_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ _12967_/A VGND VGND VPWR VPWR _12860_/A sky130_fd_sc_hd__clkbuf_1
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222_ _15209_/Q _14537_/Q _14985_/Q _15401_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14222_/X sky130_fd_sc_hd__mux4_1
X_11434_ _11434_/A VGND VGND VPWR VPWR _11434_/X sky130_fd_sc_hd__buf_1
XFILLER_138_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14153_ _14672_/Q _15248_/Q _14736_/Q _14704_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14153_/X sky130_fd_sc_hd__mux4_2
X_11365_ _11395_/A VGND VGND VPWR VPWR _11385_/A sky130_fd_sc_hd__buf_2
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13104_ _15650_/Q data_address[15] _15667_/Q VGND VGND VPWR VPWR _13104_/X sky130_fd_sc_hd__mux2_1
X_10316_ _10395_/A VGND VGND VPWR VPWR _10341_/A sky130_fd_sc_hd__buf_2
X_14084_ _15191_/Q _15159_/Q _14775_/Q _14807_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14084_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11296_ _14602_/Q _11294_/X _11174_/X _11295_/X VGND VGND VPWR VPWR _14602_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13035_ wdata[8] rdata[8] _13058_/S VGND VGND VPWR VPWR _14312_/D sky130_fd_sc_hd__mux2_4
X_10247_ _10247_/A VGND VGND VPWR VPWR _10247_/X sky130_fd_sc_hd__buf_1
XFILLER_140_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10178_ _10180_/A VGND VGND VPWR VPWR _10178_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14986_ _09786_/X _14986_/D VGND VGND VPWR VPWR _14986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13937_ _14630_/Q _14598_/Q _14566_/Q _15366_/Q _07542_/A _13950_/S1 VGND VGND VPWR
+ VPWR _13937_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13868_ _14509_/Q _14477_/Q _14445_/Q _14413_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13868_/X sky130_fd_sc_hd__mux4_1
X_12819_ _12819_/A _12927_/A VGND VGND VPWR VPWR _12967_/B sky130_fd_sc_hd__or2_1
X_15607_ _15648_/CLK _15607_/D VGND VGND VPWR VPWR pc[2] sky130_fd_sc_hd__dfxtp_1
X_13799_ _14836_/Q _14868_/Q _14900_/Q _14932_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13799_/X sky130_fd_sc_hd__mux4_2
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15538_ _15576_/CLK _15538_/D VGND VGND VPWR VPWR _15538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15469_ _15469_/CLK _15469_/D VGND VGND VPWR VPWR _15469_/Q sky130_fd_sc_hd__dfxtp_1
X_08010_ _14321_/Q VGND VGND VPWR VPWR _08011_/A sky130_fd_sc_hd__buf_1
XFILLER_118_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1 _13076_/S VGND VGND VPWR VPWR _13090_/S sky130_fd_sc_hd__buf_8
X_09961_ _09961_/A VGND VGND VPWR VPWR _09961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08912_ _08918_/A VGND VGND VPWR VPWR _08912_/X sky130_fd_sc_hd__clkbuf_1
X_09892_ _09910_/A VGND VGND VPWR VPWR _09897_/A sky130_fd_sc_hd__buf_1
XFILLER_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08843_ _08843_/A VGND VGND VPWR VPWR _08843_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08774_ _08807_/A VGND VGND VPWR VPWR _08788_/A sky130_fd_sc_hd__buf_1
XFILLER_66_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07725_ _07725_/A VGND VGND VPWR VPWR _07725_/X sky130_fd_sc_hd__buf_1
XFILLER_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07656_ _07663_/A VGND VGND VPWR VPWR _07786_/A sky130_fd_sc_hd__buf_1
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07587_ _07809_/A VGND VGND VPWR VPWR _07596_/A sky130_fd_sc_hd__buf_1
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09326_ _09335_/A VGND VGND VPWR VPWR _09326_/X sky130_fd_sc_hd__buf_1
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09257_ _09269_/A VGND VGND VPWR VPWR _09266_/A sky130_fd_sc_hd__buf_1
XFILLER_138_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08208_ _15366_/Q _08204_/X _08084_/X _08205_/X VGND VGND VPWR VPWR _15366_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09188_ _09188_/A VGND VGND VPWR VPWR _09188_/X sky130_fd_sc_hd__buf_1
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08139_ _08139_/A VGND VGND VPWR VPWR _08139_/X sky130_fd_sc_hd__clkbuf_1
X_11150_ _14640_/Q _11147_/X _11148_/X _11149_/X VGND VGND VPWR VPWR _14640_/D sky130_fd_sc_hd__a22o_1
XFILLER_107_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10101_ _14907_/Q _10097_/X _09962_/X _10098_/X VGND VGND VPWR VPWR _14907_/D sky130_fd_sc_hd__a22o_1
X_11081_ _11449_/A VGND VGND VPWR VPWR _11081_/X sky130_fd_sc_hd__buf_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10032_ _10032_/A VGND VGND VPWR VPWR _10041_/A sky130_fd_sc_hd__buf_1
XFILLER_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14840_ _10343_/X _14840_/D VGND VGND VPWR VPWR _14840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14771_ _10606_/X _14771_/D VGND VGND VPWR VPWR _14771_/Q sky130_fd_sc_hd__dfxtp_1
X_11983_ _11994_/A VGND VGND VPWR VPWR _11992_/A sky130_fd_sc_hd__buf_1
XFILLER_17_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13722_ _15227_/Q _14555_/Q _15003_/Q _15419_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13722_/X sky130_fd_sc_hd__mux4_1
X_10934_ _10956_/A VGND VGND VPWR VPWR _10941_/A sky130_fd_sc_hd__buf_1
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13653_ _14690_/Q _15266_/Q _14754_/Q _14722_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13653_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10865_ _10875_/A VGND VGND VPWR VPWR _10865_/X sky130_fd_sc_hd__buf_1
XFILLER_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12604_ _12909_/A VGND VGND VPWR VPWR _12604_/Y sky130_fd_sc_hd__inv_2
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13584_ _14126_/X _14131_/X _13648_/S VGND VGND VPWR VPWR _13584_/X sky130_fd_sc_hd__mux2_1
X_10796_ _10802_/A VGND VGND VPWR VPWR _10796_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15323_ _08393_/X _15323_/D VGND VGND VPWR VPWR _15323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12535_ _12681_/A VGND VGND VPWR VPWR _12535_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15254_ _08710_/X _15254_/D VGND VGND VPWR VPWR _15254_/Q sky130_fd_sc_hd__dfxtp_1
X_12466_ _12466_/A _12509_/B VGND VGND VPWR VPWR _12466_/Y sky130_fd_sc_hd__nor2_2
XFILLER_126_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14205_ _15115_/Q _15339_/Q _15307_/Q _15275_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14205_/X sky130_fd_sc_hd__mux4_2
X_11417_ _11424_/A VGND VGND VPWR VPWR _11422_/A sky130_fd_sc_hd__buf_1
XFILLER_126_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15185_ _08989_/X _15185_/D VGND VGND VPWR VPWR _15185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12397_ _12432_/A _12397_/B VGND VGND VPWR VPWR _12410_/B sky130_fd_sc_hd__nor2_2
XFILLER_125_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14136_ _14132_/X _14133_/X _14134_/X _14135_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14136_/X sky130_fd_sc_hd__mux4_2
X_11348_ _11368_/A VGND VGND VPWR VPWR _11353_/A sky130_fd_sc_hd__buf_2
XFILLER_126_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14067_ _14649_/Q _14617_/Q _14585_/Q _15385_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14067_/X sky130_fd_sc_hd__mux4_2
X_11279_ _14606_/Q _11273_/X _11156_/X _11274_/X VGND VGND VPWR VPWR _14606_/D sky130_fd_sc_hd__a22o_1
X_13018_ _14362_/Q VGND VGND VPWR VPWR _13018_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14969_ _09845_/X _14969_/D VGND VGND VPWR VPWR _14969_/Q sky130_fd_sc_hd__dfxtp_1
X_07510_ _07510_/A _07510_/B VGND VGND VPWR VPWR _15515_/D sky130_fd_sc_hd__nor2_1
X_08490_ _14313_/Q VGND VGND VPWR VPWR _10787_/A sky130_fd_sc_hd__buf_1
XFILLER_23_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07441_ _07442_/A _13647_/X VGND VGND VPWR VPWR _15562_/D sky130_fd_sc_hd__and2_1
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07372_ _14397_/Q VGND VGND VPWR VPWR _12571_/A sky130_fd_sc_hd__inv_2
X_09111_ _15151_/Q _09106_/X _08869_/X _09107_/X VGND VGND VPWR VPWR _15151_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09042_ _09052_/A VGND VGND VPWR VPWR _09055_/A sky130_fd_sc_hd__inv_2
XFILLER_128_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09944_ _10314_/A VGND VGND VPWR VPWR _09944_/X sky130_fd_sc_hd__buf_1
XFILLER_131_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09875_ _14961_/Q _09868_/X _09622_/X _09869_/X VGND VGND VPWR VPWR _14961_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08826_ _09196_/A VGND VGND VPWR VPWR _08826_/X sky130_fd_sc_hd__buf_1
XFILLER_58_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08757_ _08761_/A VGND VGND VPWR VPWR _08757_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07708_ _07841_/A VGND VGND VPWR VPWR _07777_/C sky130_fd_sc_hd__inv_2
X_08688_ _08692_/A VGND VGND VPWR VPWR _08688_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07639_ _07835_/A VGND VGND VPWR VPWR _07640_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10650_ _10674_/A VGND VGND VPWR VPWR _10655_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09309_ _09309_/A VGND VGND VPWR VPWR _09374_/A sky130_fd_sc_hd__buf_2
XFILLER_139_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10581_ _10583_/A VGND VGND VPWR VPWR _10581_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12320_ _12867_/A VGND VGND VPWR VPWR _12343_/A sky130_fd_sc_hd__buf_1
XFILLER_139_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12251_ _15566_/Q VGND VGND VPWR VPWR _12251_/X sky130_fd_sc_hd__buf_1
XFILLER_108_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11202_ _14627_/Q _11064_/A _11201_/X _11068_/A VGND VGND VPWR VPWR _14627_/D sky130_fd_sc_hd__a22o_1
X_12182_ _15540_/Q VGND VGND VPWR VPWR _12752_/A sky130_fd_sc_hd__buf_1
XFILLER_108_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11133_ _11147_/A VGND VGND VPWR VPWR _11133_/X sky130_fd_sc_hd__buf_1
XFILLER_89_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11064_ _11064_/A VGND VGND VPWR VPWR _11064_/X sky130_fd_sc_hd__buf_1
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10015_ _10015_/A VGND VGND VPWR VPWR _10015_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14823_ _10417_/X _14823_/D VGND VGND VPWR VPWR _14823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11966_ _11976_/A VGND VGND VPWR VPWR _11966_/X sky130_fd_sc_hd__buf_1
X_14754_ _10660_/X _14754_/D VGND VGND VPWR VPWR _14754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10917_ _14701_/Q _10914_/X _10782_/X _10916_/X VGND VGND VPWR VPWR _14701_/D sky130_fd_sc_hd__a22o_1
X_13705_ _15133_/Q _15357_/Q _15325_/Q _15293_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13705_/X sky130_fd_sc_hd__mux4_2
X_14685_ _10973_/X _14685_/D VGND VGND VPWR VPWR _14685_/Q sky130_fd_sc_hd__dfxtp_1
X_11897_ _14439_/Q _11895_/X _08079_/A _11896_/X VGND VGND VPWR VPWR _14439_/D sky130_fd_sc_hd__a22o_1
X_13636_ _14256_/X _14261_/X _13648_/S VGND VGND VPWR VPWR _13636_/X sky130_fd_sc_hd__mux2_2
X_10848_ _14720_/Q _10840_/X _10677_/X _10843_/X VGND VGND VPWR VPWR _14720_/D sky130_fd_sc_hd__a22o_1
X_13567_ _13566_/X _13080_/X _14337_/Q VGND VGND VPWR VPWR _13567_/X sky130_fd_sc_hd__mux2_1
X_10779_ _10779_/A VGND VGND VPWR VPWR _10812_/A sky130_fd_sc_hd__buf_1
XFILLER_12_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12518_ _12522_/A _12518_/B VGND VGND VPWR VPWR _12519_/B sky130_fd_sc_hd__or2_2
X_15306_ _08501_/X _15306_/D VGND VGND VPWR VPWR _15306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13498_ _13497_/X rdata[8] _13516_/S VGND VGND VPWR VPWR _13498_/X sky130_fd_sc_hd__mux2_4
X_15237_ _08768_/X _15237_/D VGND VGND VPWR VPWR _15237_/Q sky130_fd_sc_hd__dfxtp_1
X_12449_ _12593_/A _12447_/Y _12448_/X VGND VGND VPWR VPWR _12449_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15168_ _09049_/X _15168_/D VGND VGND VPWR VPWR _15168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14119_ _14836_/Q _14868_/Q _14900_/Q _14932_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14119_/X sky130_fd_sc_hd__mux4_2
X_07990_ _08038_/A VGND VGND VPWR VPWR _08023_/A sky130_fd_sc_hd__clkbuf_2
X_15099_ _09329_/X _15099_/D VGND VGND VPWR VPWR _15099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09660_ _09675_/A VGND VGND VPWR VPWR _09660_/X sky130_fd_sc_hd__buf_1
XFILLER_67_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08611_ _15282_/Q _08607_/X _08454_/X _08608_/X VGND VGND VPWR VPWR _15282_/D sky130_fd_sc_hd__a22o_1
XFILLER_94_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09591_ _09599_/A VGND VGND VPWR VPWR _09591_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08542_ _08542_/A VGND VGND VPWR VPWR _08542_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08473_ _15311_/Q _08463_/X _08472_/X _08467_/X VGND VGND VPWR VPWR _15311_/D sky130_fd_sc_hd__a22o_1
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07424_ _07424_/A _13603_/X VGND VGND VPWR VPWR _15573_/D sky130_fd_sc_hd__and2_1
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07355_ _14382_/Q VGND VGND VPWR VPWR _07506_/B sky130_fd_sc_hd__inv_2
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07286_ _07286_/A _07286_/B VGND VGND VPWR VPWR _15610_/D sky130_fd_sc_hd__nor2_1
XFILLER_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09025_ _09025_/A VGND VGND VPWR VPWR _09025_/X sky130_fd_sc_hd__buf_1
XFILLER_136_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09927_ _09927_/A VGND VGND VPWR VPWR _09927_/X sky130_fd_sc_hd__buf_1
XFILLER_77_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09858_ _09878_/A VGND VGND VPWR VPWR _09858_/X sky130_fd_sc_hd__buf_1
XFILLER_85_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08809_ _09180_/A VGND VGND VPWR VPWR _08809_/X sky130_fd_sc_hd__buf_1
X_09789_ _14986_/Q _09787_/X _09662_/X _09788_/X VGND VGND VPWR VPWR _14986_/D sky130_fd_sc_hd__a22o_1
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_103 pc[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11820_ _11820_/A VGND VGND VPWR VPWR _11839_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_114 pc[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 rdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_136 rdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_147 rdata[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_158 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11751_ _11751_/A VGND VGND VPWR VPWR _11751_/X sky130_fd_sc_hd__buf_1
XFILLER_14_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_169 wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10702_ _10702_/A VGND VGND VPWR VPWR _11463_/A sky130_fd_sc_hd__clkbuf_2
X_14470_ _11788_/X _14470_/D VGND VGND VPWR VPWR _14470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11682_ _14500_/Q _11578_/A _11567_/X _11581_/A VGND VGND VPWR VPWR _14500_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13421_ _12974_/A _12984_/X _13421_/S VGND VGND VPWR VPWR _13421_/X sky130_fd_sc_hd__mux2_1
X_10633_ _14764_/Q _10627_/X _10399_/X _10629_/X VGND VGND VPWR VPWR _14764_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13352_ _13413_/X _13411_/X _13415_/S VGND VGND VPWR VPWR _13352_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10564_ _10584_/A VGND VGND VPWR VPWR _10564_/X sky130_fd_sc_hd__buf_1
X_12303_ _12329_/A _12303_/B VGND VGND VPWR VPWR _12357_/A sky130_fd_sc_hd__nor2_4
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13283_ _12775_/X _12812_/A _13418_/S VGND VGND VPWR VPWR _13283_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10495_ _10501_/A VGND VGND VPWR VPWR _10495_/X sky130_fd_sc_hd__clkbuf_1
X_15022_ _09635_/X _15022_/D VGND VGND VPWR VPWR _15022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12234_ _12805_/A VGND VGND VPWR VPWR _12806_/A sky130_fd_sc_hd__inv_2
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12165_ _15573_/Q VGND VGND VPWR VPWR _12737_/B sky130_fd_sc_hd__inv_2
XFILLER_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11116_ _11484_/A VGND VGND VPWR VPWR _11116_/X sky130_fd_sc_hd__buf_1
XFILLER_96_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12096_ _15549_/Q VGND VGND VPWR VPWR _12626_/A sky130_fd_sc_hd__buf_1
XFILLER_110_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11047_ _11047_/A VGND VGND VPWR VPWR _11047_/X sky130_fd_sc_hd__buf_1
XFILLER_76_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14806_ _10482_/X _14806_/D VGND VGND VPWR VPWR _14806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12998_ _14342_/Q VGND VGND VPWR VPWR _12998_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14737_ _10759_/X _14737_/D VGND VGND VPWR VPWR _14737_/Q sky130_fd_sc_hd__dfxtp_1
X_11949_ _11951_/A VGND VGND VPWR VPWR _11949_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14668_ _11032_/X _14668_/D VGND VGND VPWR VPWR _14668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13619_ _13618_/X _13067_/X _14337_/Q VGND VGND VPWR VPWR _13619_/X sky130_fd_sc_hd__mux2_1
X_14599_ _11302_/X _14599_/D VGND VGND VPWR VPWR _14599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07140_ _13104_/X VGND VGND VPWR VPWR _07272_/B sky130_fd_sc_hd__inv_2
XFILLER_118_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07973_ _07973_/A VGND VGND VPWR VPWR _07973_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09712_ _09722_/A VGND VGND VPWR VPWR _09712_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09643_ _10394_/A VGND VGND VPWR VPWR _09643_/X sky130_fd_sc_hd__buf_1
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09574_ _10336_/A VGND VGND VPWR VPWR _09574_/X sky130_fd_sc_hd__buf_1
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08525_ _15303_/Q _08520_/X _08523_/X _08524_/X VGND VGND VPWR VPWR _15303_/D sky130_fd_sc_hd__a22o_1
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ _08474_/A VGND VGND VPWR VPWR _08469_/A sky130_fd_sc_hd__buf_1
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07407_ _07420_/A VGND VGND VPWR VPWR _07416_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08387_ _08405_/A VGND VGND VPWR VPWR _08387_/X sky130_fd_sc_hd__buf_1
X_07338_ _07338_/A VGND VGND VPWR VPWR _07354_/A sky130_fd_sc_hd__buf_1
XFILLER_109_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07269_ _07269_/A _07269_/B VGND VGND VPWR VPWR _15622_/D sky130_fd_sc_hd__nor2_1
X_09008_ _09026_/A VGND VGND VPWR VPWR _09008_/X sky130_fd_sc_hd__buf_1
X_10280_ _10280_/A VGND VGND VPWR VPWR _10280_/X sky130_fd_sc_hd__buf_1
XFILLER_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13970_ _14947_/Q _15043_/Q _15011_/Q _15075_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13970_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12921_ _12315_/A _12854_/X _12852_/X _12838_/A VGND VGND VPWR VPWR _12924_/B sky130_fd_sc_hd__o22a_1
XFILLER_86_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15640_ _15648_/CLK _15640_/D VGND VGND VPWR VPWR _15640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12852_ _12852_/A VGND VGND VPWR VPWR _12852_/X sky130_fd_sc_hd__buf_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11803_ _11803_/A VGND VGND VPWR VPWR _11803_/X sky130_fd_sc_hd__buf_1
X_15571_ _15576_/CLK _15571_/D VGND VGND VPWR VPWR _15571_/Q sky130_fd_sc_hd__dfxtp_1
X_12783_ _12783_/A VGND VGND VPWR VPWR _12810_/A sky130_fd_sc_hd__buf_1
XFILLER_42_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_53_clk _14315_/CLK VGND VGND VPWR VPWR _15663_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11734_ _11765_/A VGND VGND VPWR VPWR _11753_/A sky130_fd_sc_hd__clkbuf_2
X_14522_ _11608_/X _14522_/D VGND VGND VPWR VPWR _14522_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14453_ _11848_/X _14453_/D VGND VGND VPWR VPWR _14453_/Q sky130_fd_sc_hd__dfxtp_1
X_11665_ _11674_/A VGND VGND VPWR VPWR _11665_/X sky130_fd_sc_hd__buf_1
XFILLER_30_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _12611_/X _12610_/X _13418_/S VGND VGND VPWR VPWR _13404_/X sky130_fd_sc_hd__mux2_1
X_10616_ _10616_/A VGND VGND VPWR VPWR _10616_/X sky130_fd_sc_hd__buf_1
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ _14393_/CLK instruction[13] VGND VGND VPWR VPWR _14384_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11596_ _11598_/A VGND VGND VPWR VPWR _11596_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13335_ _13377_/X _13374_/X _13415_/S VGND VGND VPWR VPWR _13335_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10547_ _10547_/A VGND VGND VPWR VPWR _10547_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13266_ _13334_/X _13331_/X _13393_/S VGND VGND VPWR VPWR _13266_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10478_ _14808_/Q _10474_/X _10344_/X _10475_/X VGND VGND VPWR VPWR _14808_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12217_ _15531_/Q VGND VGND VPWR VPWR _12862_/A sky130_fd_sc_hd__inv_2
X_15005_ _09722_/X _15005_/D VGND VGND VPWR VPWR _15005_/Q sky130_fd_sc_hd__dfxtp_1
X_13197_ _12329_/X _12590_/X _13418_/S VGND VGND VPWR VPWR _13197_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12148_ _12148_/A VGND VGND VPWR VPWR _12148_/X sky130_fd_sc_hd__buf_1
XFILLER_96_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12079_ _15584_/Q VGND VGND VPWR VPWR _12079_/X sky130_fd_sc_hd__buf_1
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk _14315_/CLK VGND VGND VPWR VPWR _15599_/CLK sky130_fd_sc_hd__clkbuf_16
X_08310_ _08319_/A VGND VGND VPWR VPWR _08315_/A sky130_fd_sc_hd__buf_1
X_09290_ _09290_/A VGND VGND VPWR VPWR _09290_/X sky130_fd_sc_hd__buf_1
X_08241_ _08261_/A VGND VGND VPWR VPWR _08241_/X sky130_fd_sc_hd__buf_1
XANTENNA_14 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 data_address[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08172_ _08178_/A VGND VGND VPWR VPWR _08172_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_58 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 pc[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07123_ _07123_/A VGND VGND VPWR VPWR _13152_/S sky130_fd_sc_hd__inv_16
XFILLER_146_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07956_ _07956_/A VGND VGND VPWR VPWR _07956_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07887_ _07731_/X _07885_/Y _07874_/X _07820_/A _07886_/Y VGND VGND VPWR VPWR _15436_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09626_ _10765_/A VGND VGND VPWR VPWR _10379_/A sky130_fd_sc_hd__buf_1
XFILLER_83_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09557_ _09567_/A VGND VGND VPWR VPWR _09557_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_clk _14397_/CLK VGND VGND VPWR VPWR _15576_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08508_ _08508_/A VGND VGND VPWR VPWR _08508_/X sky130_fd_sc_hd__clkbuf_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09488_ _09506_/A VGND VGND VPWR VPWR _09488_/X sky130_fd_sc_hd__buf_1
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ _08451_/A VGND VGND VPWR VPWR _08439_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11450_ _11450_/A VGND VGND VPWR VPWR _11529_/A sky130_fd_sc_hd__clkbuf_4
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10401_ _10413_/A VGND VGND VPWR VPWR _10410_/A sky130_fd_sc_hd__buf_1
XFILLER_137_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11381_ _11383_/A VGND VGND VPWR VPWR _11381_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13120_ _15666_/Q data_address[31] _15667_/Q VGND VGND VPWR VPWR _13120_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10332_ _10332_/A VGND VGND VPWR VPWR _10332_/X sky130_fd_sc_hd__buf_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13051_ wdata[24] rdata[24] _13057_/S VGND VGND VPWR VPWR _14328_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10263_ _14860_/Q _10257_/X _10030_/X _10259_/X VGND VGND VPWR VPWR _14860_/D sky130_fd_sc_hd__a22o_1
XFILLER_127_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12002_ _14408_/Q _11996_/X _08074_/A _11997_/X VGND VGND VPWR VPWR _14408_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10194_ _10194_/A VGND VGND VPWR VPWR _10256_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13953_ _14660_/Q _15236_/Q _14724_/Q _14692_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13953_/X sky130_fd_sc_hd__mux4_2
XFILLER_47_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12904_ _12904_/A _12904_/B _12904_/C _12904_/D VGND VGND VPWR VPWR _12905_/C sky130_fd_sc_hd__or4_4
XFILLER_62_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13884_ _15179_/Q _15147_/Q _14763_/Q _14795_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13884_/X sky130_fd_sc_hd__mux4_2
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15623_ _15654_/CLK _15623_/D VGND VGND VPWR VPWR pc[18] sky130_fd_sc_hd__dfxtp_1
X_12835_ _13296_/X VGND VGND VPWR VPWR _12835_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_26_clk _14397_/CLK VGND VGND VPWR VPWR _14392_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15554_ _15589_/CLK _15554_/D VGND VGND VPWR VPWR _15554_/Q sky130_fd_sc_hd__dfxtp_1
X_12766_ _12762_/X _12763_/X _12715_/X VGND VGND VPWR VPWR _12766_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14505_ _11667_/X _14505_/D VGND VGND VPWR VPWR _14505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11717_ _11721_/A VGND VGND VPWR VPWR _11717_/X sky130_fd_sc_hd__clkbuf_1
X_15485_ _15510_/CLK _15485_/D VGND VGND VPWR VPWR wdata[11] sky130_fd_sc_hd__dfxtp_4
X_12697_ _12740_/A VGND VGND VPWR VPWR _12826_/A sky130_fd_sc_hd__buf_1
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _14510_/Q _11642_/X _11523_/X _11643_/X VGND VGND VPWR VPWR _14510_/D sky130_fd_sc_hd__a22o_1
X_14436_ _11903_/X _14436_/D VGND VGND VPWR VPWR _14436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14367_ _14392_/CLK pc[28] VGND VGND VPWR VPWR _14367_/Q sky130_fd_sc_hd__dfxtp_1
X_11579_ _11589_/A VGND VGND VPWR VPWR _11592_/A sky130_fd_sc_hd__inv_2
X_13318_ _13317_/X _13319_/X _15565_/Q VGND VGND VPWR VPWR _13318_/X sky130_fd_sc_hd__mux2_1
X_14298_ _15510_/CLK _15465_/Q VGND VGND VPWR VPWR _14298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13249_ _13248_/X _12489_/X _15565_/Q VGND VGND VPWR VPWR _13249_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07810_ _07869_/A VGND VGND VPWR VPWR _07810_/X sky130_fd_sc_hd__buf_1
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08790_ _15233_/Q _08782_/X _08789_/X _08786_/X VGND VGND VPWR VPWR _15233_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07741_ _07739_/X _07740_/X _07739_/X _07740_/X VGND VGND VPWR VPWR _07891_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_38_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07672_ _07670_/X _07671_/X _07670_/X _13126_/X VGND VGND VPWR VPWR _07803_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09411_ _09423_/A VGND VGND VPWR VPWR _09426_/A sky130_fd_sc_hd__inv_2
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_clk _14397_/CLK VGND VGND VPWR VPWR _15505_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09342_ _09342_/A VGND VGND VPWR VPWR _09351_/A sky130_fd_sc_hd__buf_1
XFILLER_80_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09273_ _09278_/A VGND VGND VPWR VPWR _09273_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08224_ _08660_/A VGND VGND VPWR VPWR _11686_/A sky130_fd_sc_hd__buf_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08155_ _08174_/A VGND VGND VPWR VPWR _08155_/X sky130_fd_sc_hd__buf_1
X_07106_ _07383_/A VGND VGND VPWR VPWR _07642_/A sky130_fd_sc_hd__buf_1
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08086_ _08191_/A VGND VGND VPWR VPWR _08161_/A sky130_fd_sc_hd__buf_1
XFILLER_134_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08988_ _15186_/Q _08984_/X _08856_/X _08985_/X VGND VGND VPWR VPWR _15186_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07939_ _08191_/A VGND VGND VPWR VPWR _08038_/A sky130_fd_sc_hd__buf_2
XFILLER_44_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10950_ _10962_/A VGND VGND VPWR VPWR _10951_/A sky130_fd_sc_hd__buf_1
XFILLER_44_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09609_ _09615_/A VGND VGND VPWR VPWR _09609_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10881_ _10892_/A VGND VGND VPWR VPWR _10890_/A sky130_fd_sc_hd__buf_1
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12620_ _12620_/A VGND VGND VPWR VPWR _12620_/X sky130_fd_sc_hd__buf_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ _12551_/A _15464_/Q VGND VGND VPWR VPWR _12551_/Y sky130_fd_sc_hd__nor2_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11502_ _11502_/A VGND VGND VPWR VPWR _11502_/X sky130_fd_sc_hd__buf_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _12460_/X _12469_/Y _12477_/Y _12481_/X VGND VGND VPWR VPWR _12482_/Y sky130_fd_sc_hd__o211ai_2
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15270_ _08650_/X _15270_/D VGND VGND VPWR VPWR _15270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11433_ _11450_/A VGND VGND VPWR VPWR _11434_/A sky130_fd_sc_hd__buf_1
X_14221_ _14217_/X _14218_/X _14219_/X _14220_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14221_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14152_ _15216_/Q _14544_/Q _14992_/Q _15408_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14152_/X sky130_fd_sc_hd__mux4_1
X_11364_ _11384_/A VGND VGND VPWR VPWR _11364_/X sky130_fd_sc_hd__buf_1
XFILLER_152_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13103_ _15649_/Q data_address[14] _15667_/Q VGND VGND VPWR VPWR _13103_/X sky130_fd_sc_hd__mux2_1
X_10315_ _10315_/A VGND VGND VPWR VPWR _10395_/A sky130_fd_sc_hd__buf_2
X_14083_ _14679_/Q _15255_/Q _14743_/Q _14711_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14083_/X sky130_fd_sc_hd__mux4_2
X_11295_ _11304_/A VGND VGND VPWR VPWR _11295_/X sky130_fd_sc_hd__buf_1
XFILLER_125_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13034_ wdata[7] rdata[7] _13058_/S VGND VGND VPWR VPWR _14311_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10246_ _10246_/A VGND VGND VPWR VPWR _10246_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10177_ _14884_/Q _10071_/A _10062_/X _10074_/A VGND VGND VPWR VPWR _14884_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14985_ _09790_/X _14985_/D VGND VGND VPWR VPWR _14985_/Q sky130_fd_sc_hd__dfxtp_1
X_13936_ _13932_/X _13933_/X _13934_/X _13935_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13936_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13867_ _14637_/Q _14605_/Q _14573_/Q _15373_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13867_/X sky130_fd_sc_hd__mux4_2
X_15606_ _15669_/CLK _15606_/D VGND VGND VPWR VPWR pc[1] sky130_fd_sc_hd__dfxtp_1
X_12818_ _12926_/A _12926_/B VGND VGND VPWR VPWR _12927_/A sky130_fd_sc_hd__nand2_1
XFILLER_90_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13798_ _14516_/Q _14484_/Q _14452_/Q _14420_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13798_/X sky130_fd_sc_hd__mux4_1
X_15537_ _15576_/CLK _15537_/D VGND VGND VPWR VPWR _15537_/Q sky130_fd_sc_hd__dfxtp_1
X_12749_ _12749_/A _12749_/B VGND VGND VPWR VPWR _12750_/B sky130_fd_sc_hd__nand2_2
X_15468_ _15469_/CLK _15468_/D VGND VGND VPWR VPWR _15468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14419_ _11965_/X _14419_/D VGND VGND VPWR VPWR _14419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15399_ _08076_/X _15399_/D VGND VGND VPWR VPWR _15399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater2 _14338_/Q VGND VGND VPWR VPWR _13516_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_116_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09960_ _14940_/Q _09957_/X _09958_/X _09959_/X VGND VGND VPWR VPWR _14940_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_6_clk clkbuf_opt_4_clk/X VGND VGND VPWR VPWR _14399_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08911_ _08921_/A VGND VGND VPWR VPWR _08918_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09891_ _09917_/A VGND VGND VPWR VPWR _09910_/A sky130_fd_sc_hd__buf_1
XFILLER_112_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08842_ _15222_/Q _08838_/X _08839_/X _08841_/X VGND VGND VPWR VPWR _15222_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08773_ _08858_/A VGND VGND VPWR VPWR _08807_/A sky130_fd_sc_hd__buf_1
X_07724_ _15603_/Q VGND VGND VPWR VPWR _07725_/A sky130_fd_sc_hd__inv_2
XFILLER_38_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07655_ _07655_/A VGND VGND VPWR VPWR _07663_/A sky130_fd_sc_hd__buf_1
XFILLER_80_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07586_ _07586_/A VGND VGND VPWR VPWR _07809_/A sky130_fd_sc_hd__buf_1
XFILLER_41_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09325_ _09331_/A VGND VGND VPWR VPWR _09325_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09256_ _15116_/Q _09249_/X _09255_/X _09252_/X VGND VGND VPWR VPWR _15116_/D sky130_fd_sc_hd__a22o_1
X_08207_ _08209_/A VGND VGND VPWR VPWR _08207_/X sky130_fd_sc_hd__clkbuf_1
X_09187_ _09187_/A VGND VGND VPWR VPWR _09187_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08138_ _15387_/Q _08134_/X _07973_/X _08135_/X VGND VGND VPWR VPWR _15387_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08069_ _08069_/A VGND VGND VPWR VPWR _08069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10100_ _10102_/A VGND VGND VPWR VPWR _10100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11080_ _11107_/A VGND VGND VPWR VPWR _11080_/X sky130_fd_sc_hd__buf_1
XFILLER_49_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10031_ _14924_/Q _10024_/X _10030_/X _10027_/X VGND VGND VPWR VPWR _14924_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14770_ _10611_/X _14770_/D VGND VGND VPWR VPWR _14770_/Q sky130_fd_sc_hd__dfxtp_1
X_11982_ _14414_/Q _11976_/X _08042_/A _11977_/X VGND VGND VPWR VPWR _14414_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13721_ _13717_/X _13718_/X _13719_/X _13720_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13721_/X sky130_fd_sc_hd__mux4_1
X_10933_ _10999_/A VGND VGND VPWR VPWR _10956_/A sky130_fd_sc_hd__buf_2
XFILLER_56_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10864_ _10874_/A VGND VGND VPWR VPWR _10864_/X sky130_fd_sc_hd__buf_1
X_13652_ _15234_/Q _14562_/Q _15010_/Q _15426_/Q _13740_/S0 _07541_/A VGND VGND VPWR
+ VPWR _13652_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12603_ _12599_/X _12577_/X _12065_/X _12602_/X VGND VGND VPWR VPWR _12909_/A sky130_fd_sc_hd__o22a_1
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10795_ _14731_/Q _10780_/X _10794_/X _10784_/X VGND VGND VPWR VPWR _14731_/D sky130_fd_sc_hd__a22o_1
X_13583_ _13582_/X _13076_/X _14337_/Q VGND VGND VPWR VPWR _13583_/X sky130_fd_sc_hd__mux2_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15322_ _08399_/X _15322_/D VGND VGND VPWR VPWR _15322_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12534_ _12534_/A VGND VGND VPWR VPWR _12534_/Y sky130_fd_sc_hd__inv_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15253_ _08718_/X _15253_/D VGND VGND VPWR VPWR _15253_/Q sky130_fd_sc_hd__dfxtp_1
X_12465_ _12463_/X _12347_/X _12473_/A _12505_/A VGND VGND VPWR VPWR _12509_/B sky130_fd_sc_hd__o22a_2
XFILLER_138_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14204_ _15179_/Q _15147_/Q _14763_/Q _14795_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14204_/X sky130_fd_sc_hd__mux4_2
X_11416_ _14567_/Q _11414_/X _11187_/X _11415_/X VGND VGND VPWR VPWR _14567_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15184_ _08992_/X _15184_/D VGND VGND VPWR VPWR _15184_/Q sky130_fd_sc_hd__dfxtp_1
X_12396_ _12355_/Y _12357_/X _12395_/Y VGND VGND VPWR VPWR _12397_/B sky130_fd_sc_hd__o21ai_2
XFILLER_153_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14135_ _15122_/Q _15346_/Q _15314_/Q _15282_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14135_/X sky130_fd_sc_hd__mux4_2
X_11347_ _11407_/A VGND VGND VPWR VPWR _11368_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14066_ _14062_/X _14063_/X _14064_/X _14065_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14066_/X sky130_fd_sc_hd__mux4_2
X_11278_ _11278_/A VGND VGND VPWR VPWR _11278_/X sky130_fd_sc_hd__clkbuf_1
X_13017_ _14361_/Q VGND VGND VPWR VPWR _13017_/Y sky130_fd_sc_hd__inv_2
X_10229_ _10248_/A VGND VGND VPWR VPWR _10229_/X sky130_fd_sc_hd__buf_1
XFILLER_67_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14968_ _09850_/X _14968_/D VGND VGND VPWR VPWR _14968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13919_ _14824_/Q _14856_/Q _14888_/Q _14920_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13919_/X sky130_fd_sc_hd__mux4_2
X_14899_ _10126_/X _14899_/D VGND VGND VPWR VPWR _14899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07440_ _07442_/A _13643_/X VGND VGND VPWR VPWR _15563_/D sky130_fd_sc_hd__and2_1
XFILLER_50_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07371_ _14380_/Q VGND VGND VPWR VPWR _07509_/B sky130_fd_sc_hd__inv_2
XFILLER_15_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09110_ _09114_/A VGND VGND VPWR VPWR _09110_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09041_ _09041_/A VGND VGND VPWR VPWR _09041_/X sky130_fd_sc_hd__buf_1
XFILLER_136_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09943_ _09972_/A VGND VGND VPWR VPWR _09943_/X sky130_fd_sc_hd__buf_1
XFILLER_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09874_ _09876_/A VGND VGND VPWR VPWR _09874_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08825_ _08825_/A VGND VGND VPWR VPWR _08825_/X sky130_fd_sc_hd__buf_1
XFILLER_39_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08756_ _08765_/A VGND VGND VPWR VPWR _08761_/A sky130_fd_sc_hd__buf_1
XFILLER_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07707_ _07706_/X _07683_/X _07706_/X _13134_/X VGND VGND VPWR VPWR _07841_/A sky130_fd_sc_hd__a2bb2o_1
X_08687_ _08705_/A VGND VGND VPWR VPWR _08692_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07638_ _07638_/A _15510_/Q VGND VGND VPWR VPWR _15462_/D sky130_fd_sc_hd__and2_1
XFILLER_81_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07569_ _07569_/A VGND VGND VPWR VPWR _07572_/A sky130_fd_sc_hd__clkbuf_2
X_09308_ _09318_/A VGND VGND VPWR VPWR _09308_/X sky130_fd_sc_hd__clkbuf_1
X_10580_ _14779_/Q _10575_/X _10332_/X _10576_/X VGND VGND VPWR VPWR _14779_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09239_ _09239_/A VGND VGND VPWR VPWR _09239_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12250_ _12254_/A VGND VGND VPWR VPWR _12836_/A sky130_fd_sc_hd__buf_1
XFILLER_119_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11201_ _11570_/A VGND VGND VPWR VPWR _11201_/X sky130_fd_sc_hd__buf_1
X_12181_ _12179_/X _12102_/A _12755_/A _12106_/A VGND VGND VPWR VPWR _12183_/A sky130_fd_sc_hd__o22a_1
XFILLER_134_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11132_ _11137_/A VGND VGND VPWR VPWR _11132_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11063_ _11078_/A VGND VGND VPWR VPWR _11064_/A sky130_fd_sc_hd__buf_1
XFILLER_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10014_ _14928_/Q _10011_/X _10012_/X _10013_/X VGND VGND VPWR VPWR _14928_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14822_ _10422_/X _14822_/D VGND VGND VPWR VPWR _14822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14753_ _10670_/X _14753_/D VGND VGND VPWR VPWR _14753_/Q sky130_fd_sc_hd__dfxtp_1
X_11965_ _11971_/A VGND VGND VPWR VPWR _11965_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13704_ _15197_/Q _15165_/Q _14781_/Q _14813_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13704_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10916_ _10937_/A VGND VGND VPWR VPWR _10916_/X sky130_fd_sc_hd__buf_1
X_14684_ _10975_/X _14684_/D VGND VGND VPWR VPWR _14684_/Q sky130_fd_sc_hd__dfxtp_1
X_11896_ _11896_/A VGND VGND VPWR VPWR _11896_/X sky130_fd_sc_hd__buf_1
XFILLER_32_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13635_ _13634_/X _13063_/X _14337_/Q VGND VGND VPWR VPWR _13635_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10847_ _10847_/A VGND VGND VPWR VPWR _10847_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13566_ _13565_/X _14325_/D _15506_/Q VGND VGND VPWR VPWR _13566_/X sky130_fd_sc_hd__mux2_2
XFILLER_13_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10778_ _10786_/A VGND VGND VPWR VPWR _10778_/X sky130_fd_sc_hd__clkbuf_1
X_15305_ _08508_/X _15305_/D VGND VGND VPWR VPWR _15305_/Q sky130_fd_sc_hd__dfxtp_1
X_12517_ _15561_/Q VGND VGND VPWR VPWR _12518_/B sky130_fd_sc_hd__buf_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13497_ _13886_/X _13891_/X _13521_/S VGND VGND VPWR VPWR _13497_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15236_ _08770_/X _15236_/D VGND VGND VPWR VPWR _15236_/Q sky130_fd_sc_hd__dfxtp_1
X_12448_ _12448_/A VGND VGND VPWR VPWR _12448_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15167_ _09051_/X _15167_/D VGND VGND VPWR VPWR _15167_/Q sky130_fd_sc_hd__dfxtp_1
X_12379_ _12379_/A _12379_/B VGND VGND VPWR VPWR _12379_/Y sky130_fd_sc_hd__nor2_2
XFILLER_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14118_ _14516_/Q _14484_/Q _14452_/Q _14420_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14118_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15098_ _09331_/X _15098_/D VGND VGND VPWR VPWR _15098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14049_ _14843_/Q _14875_/Q _14907_/Q _14939_/Q _14395_/Q _14060_/S1 VGND VGND VPWR
+ VPWR _14049_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08610_ _08612_/A VGND VGND VPWR VPWR _08610_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09590_ _15031_/Q _09577_/X _09589_/X _09580_/X VGND VGND VPWR VPWR _15031_/D sky130_fd_sc_hd__a22o_1
XFILLER_94_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08541_ _15300_/Q _08344_/A _08540_/X _08350_/A VGND VGND VPWR VPWR _15300_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08472_ _09240_/A VGND VGND VPWR VPWR _08472_/X sky130_fd_sc_hd__buf_1
XFILLER_63_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07423_ _07424_/A _13599_/X VGND VGND VPWR VPWR _15574_/D sky130_fd_sc_hd__and2_1
XFILLER_149_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07354_ _07354_/A VGND VGND VPWR VPWR _07354_/X sky130_fd_sc_hd__buf_1
XFILLER_31_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07285_ _07286_/A _07285_/B VGND VGND VPWR VPWR _15611_/D sky130_fd_sc_hd__nor2_1
XFILLER_109_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09024_ _09030_/A VGND VGND VPWR VPWR _09024_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09926_ _09941_/A VGND VGND VPWR VPWR _09927_/A sky130_fd_sc_hd__buf_1
XFILLER_86_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09857_ _09888_/A VGND VGND VPWR VPWR _09878_/A sky130_fd_sc_hd__buf_2
XFILLER_86_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08808_ _08816_/A VGND VGND VPWR VPWR _08808_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09788_ _09798_/A VGND VGND VPWR VPWR _09788_/X sky130_fd_sc_hd__buf_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_104 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08739_ _15246_/Q _08732_/X _08478_/X _08733_/X VGND VGND VPWR VPWR _15246_/D sky130_fd_sc_hd__a22o_1
XFILLER_73_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_115 pc[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_126 rdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_137 rdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_148 rdata[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11750_ _14481_/Q _11743_/X _11510_/X _11744_/X VGND VGND VPWR VPWR _14481_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_159 wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10701_ _10716_/A VGND VGND VPWR VPWR _10701_/X sky130_fd_sc_hd__buf_1
XFILLER_14_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11681_ _11685_/A VGND VGND VPWR VPWR _11681_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13420_ _12982_/Y _12980_/X _13420_/S VGND VGND VPWR VPWR _13420_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10632_ _10636_/A VGND VGND VPWR VPWR _10632_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13351_ _13410_/X _13407_/X _13415_/S VGND VGND VPWR VPWR _13351_/X sky130_fd_sc_hd__mux2_1
X_10563_ _10626_/A VGND VGND VPWR VPWR _10584_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12302_ _12021_/X _12298_/X _12330_/A _12437_/A VGND VGND VPWR VPWR _12303_/B sky130_fd_sc_hd__o22a_1
X_13282_ _13283_/X _13297_/X _13415_/S VGND VGND VPWR VPWR _13282_/X sky130_fd_sc_hd__mux2_1
X_10494_ _10512_/A VGND VGND VPWR VPWR _10501_/A sky130_fd_sc_hd__buf_1
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15021_ _09639_/X _15021_/D VGND VGND VPWR VPWR _15021_/Q sky130_fd_sc_hd__dfxtp_1
X_12233_ _15536_/Q VGND VGND VPWR VPWR _12805_/A sky130_fd_sc_hd__buf_1
XFILLER_123_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12164_ _12164_/A VGND VGND VPWR VPWR _12164_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11115_ _11125_/A VGND VGND VPWR VPWR _11115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12095_ _12091_/X _12092_/X _12627_/A _12094_/X VGND VGND VPWR VPWR _12097_/A sky130_fd_sc_hd__o22a_1
XFILLER_68_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11046_ _11046_/A VGND VGND VPWR VPWR _11046_/X sky130_fd_sc_hd__buf_1
XFILLER_37_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14805_ _10488_/X _14805_/D VGND VGND VPWR VPWR _14805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12997_ _14341_/Q VGND VGND VPWR VPWR _12997_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14736_ _10763_/X _14736_/D VGND VGND VPWR VPWR _14736_/Q sky130_fd_sc_hd__dfxtp_1
X_11948_ _14425_/Q _11946_/X _07983_/A _11947_/X VGND VGND VPWR VPWR _14425_/D sky130_fd_sc_hd__a22o_1
XFILLER_72_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14667_ _11034_/X _14667_/D VGND VGND VPWR VPWR _14667_/Q sky130_fd_sc_hd__dfxtp_1
X_11879_ _11879_/A VGND VGND VPWR VPWR _11879_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13618_ _13617_/X _14312_/D _15506_/Q VGND VGND VPWR VPWR _13618_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14598_ _11306_/X _14598_/D VGND VGND VPWR VPWR _14598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13549_ _13548_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13549_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15219_ _08850_/X _15219_/D VGND VGND VPWR VPWR _15219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07972_ _14328_/Q VGND VGND VPWR VPWR _07973_/A sky130_fd_sc_hd__buf_1
X_09711_ _09724_/A VGND VGND VPWR VPWR _09722_/A sky130_fd_sc_hd__buf_1
XFILLER_68_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09642_ _10781_/A VGND VGND VPWR VPWR _10394_/A sky130_fd_sc_hd__buf_1
XFILLER_55_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09573_ _10712_/A VGND VGND VPWR VPWR _10336_/A sky130_fd_sc_hd__buf_1
XFILLER_36_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08524_ _08524_/A VGND VGND VPWR VPWR _08524_/X sky130_fd_sc_hd__buf_1
XFILLER_36_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08455_ _15314_/Q _08445_/X _08454_/X _08449_/X VGND VGND VPWR VPWR _15314_/D sky130_fd_sc_hd__a22o_1
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07406_ _07406_/A _13555_/X VGND VGND VPWR VPWR _15585_/D sky130_fd_sc_hd__and2_1
X_08386_ _08393_/A VGND VGND VPWR VPWR _08386_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07337_ _07337_/A _07337_/B VGND VGND VPWR VPWR _15601_/D sky130_fd_sc_hd__nor2_1
X_07268_ _07269_/A _07268_/B VGND VGND VPWR VPWR _15623_/D sky130_fd_sc_hd__nor2_1
X_09007_ _09007_/A VGND VGND VPWR VPWR _09026_/A sky130_fd_sc_hd__clkbuf_2
X_07199_ _13114_/X _07197_/Y _07198_/X _07175_/B VGND VGND VPWR VPWR _15660_/D sky130_fd_sc_hd__o211a_1
XFILLER_105_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09909_ _14951_/Q _09907_/X _09677_/X _09908_/X VGND VGND VPWR VPWR _14951_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12920_ _12842_/X _12251_/X _12254_/A _12843_/A VGND VGND VPWR VPWR _12924_/A sky130_fd_sc_hd__o22a_1
XFILLER_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12851_ _12851_/A VGND VGND VPWR VPWR _12851_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11802_ _11814_/A VGND VGND VPWR VPWR _11803_/A sky130_fd_sc_hd__buf_1
X_15570_ _15576_/CLK _15570_/D VGND VGND VPWR VPWR _15570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12782_ _12782_/A VGND VGND VPWR VPWR _12782_/X sky130_fd_sc_hd__buf_1
XFILLER_54_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14521_ _11611_/X _14521_/D VGND VGND VPWR VPWR _14521_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11733_ _11752_/A VGND VGND VPWR VPWR _11733_/X sky130_fd_sc_hd__buf_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14452_ _11853_/X _14452_/D VGND VGND VPWR VPWR _14452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11664_ _11673_/A VGND VGND VPWR VPWR _11664_/X sky130_fd_sc_hd__buf_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _12577_/X _12590_/X _13418_/S VGND VGND VPWR VPWR _13403_/X sky130_fd_sc_hd__mux2_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10615_ _10615_/A VGND VGND VPWR VPWR _10615_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14383_ _14395_/CLK instruction[12] VGND VGND VPWR VPWR _14383_/Q sky130_fd_sc_hd__dfxtp_4
X_11595_ _14527_/Q _11591_/X _11449_/X _11594_/X VGND VGND VPWR VPWR _14527_/D sky130_fd_sc_hd__a22o_1
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _13336_/X _13335_/X _13408_/S VGND VGND VPWR VPWR _13334_/X sky130_fd_sc_hd__mux2_1
X_10546_ _14787_/Q _10440_/A _10434_/X _10443_/A VGND VGND VPWR VPWR _14787_/D sky130_fd_sc_hd__a22o_1
X_13265_ _12758_/A _12762_/X _15561_/Q VGND VGND VPWR VPWR _13265_/X sky130_fd_sc_hd__mux2_1
X_10477_ _10479_/A VGND VGND VPWR VPWR _10477_/X sky130_fd_sc_hd__clkbuf_1
X_15004_ _09725_/X _15004_/D VGND VGND VPWR VPWR _15004_/Q sky130_fd_sc_hd__dfxtp_1
X_12216_ _12211_/X _12230_/B _12215_/Y VGND VGND VPWR VPWR _12216_/Y sky130_fd_sc_hd__a21oi_4
X_13196_ _13197_/X _13207_/X _13415_/S VGND VGND VPWR VPWR _13196_/X sky130_fd_sc_hd__mux2_1
X_12147_ _15576_/Q VGND VGND VPWR VPWR _12694_/A sky130_fd_sc_hd__inv_2
XFILLER_151_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12078_ _15552_/Q VGND VGND VPWR VPWR _12588_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11029_ _11140_/A VGND VGND VPWR VPWR _11101_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14719_ _10850_/X _14719_/D VGND VGND VPWR VPWR _14719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08240_ _08305_/A VGND VGND VPWR VPWR _08261_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_15 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 data_address[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08171_ _08180_/A VGND VGND VPWR VPWR _08178_/A sky130_fd_sc_hd__buf_1
XANTENNA_48 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 pc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07122_ _07634_/B _12030_/C _15511_/Q _12040_/B VGND VGND VPWR VPWR _07123_/A sky130_fd_sc_hd__or4_4
XFILLER_127_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07955_ _15423_/Q _07949_/X _07951_/X _07954_/X VGND VGND VPWR VPWR _15423_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07886_ _07731_/X _07885_/Y _07874_/X VGND VGND VPWR VPWR _07886_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09625_ _09625_/A VGND VGND VPWR VPWR _09625_/X sky130_fd_sc_hd__buf_1
XFILLER_44_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09556_ _09586_/A VGND VGND VPWR VPWR _09567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08507_ _15306_/Q _08502_/X _08505_/X _08506_/X VGND VGND VPWR VPWR _15306_/D sky130_fd_sc_hd__a22o_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09487_ _09487_/A VGND VGND VPWR VPWR _09506_/A sky130_fd_sc_hd__buf_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08438_ _08474_/A VGND VGND VPWR VPWR _08451_/A sky130_fd_sc_hd__buf_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08369_ _09170_/A VGND VGND VPWR VPWR _08369_/X sky130_fd_sc_hd__buf_1
X_10400_ _14828_/Q _10393_/X _10399_/X _10396_/X VGND VGND VPWR VPWR _14828_/D sky130_fd_sc_hd__a22o_1
X_11380_ _14578_/Q _11374_/X _11138_/X _11375_/X VGND VGND VPWR VPWR _14578_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10331_ _10331_/A VGND VGND VPWR VPWR _10331_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13050_ wdata[23] rdata[23] _13057_/S VGND VGND VPWR VPWR _14327_/D sky130_fd_sc_hd__mux2_1
X_10262_ _10266_/A VGND VGND VPWR VPWR _10262_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12001_ _12001_/A VGND VGND VPWR VPWR _12001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10193_ _10193_/A VGND VGND VPWR VPWR _10193_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13952_ _15204_/Q _14532_/Q _14980_/Q _15396_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13952_/X sky130_fd_sc_hd__mux4_2
XFILLER_143_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12903_ _12480_/A _12470_/X _12905_/B _12901_/X _12902_/X VGND VGND VPWR VPWR _12903_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_47_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13883_ _14667_/Q _15243_/Q _14731_/Q _14699_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13883_/X sky130_fd_sc_hd__mux4_2
XFILLER_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15622_ _15652_/CLK _15622_/D VGND VGND VPWR VPWR pc[17] sky130_fd_sc_hd__dfxtp_4
X_12834_ _12821_/X _12824_/X _12827_/X _12832_/Y _12833_/Y VGND VGND VPWR VPWR _12834_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_61_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15553_ _15590_/CLK _15553_/D VGND VGND VPWR VPWR _15553_/Q sky130_fd_sc_hd__dfxtp_1
X_12765_ _15539_/Q VGND VGND VPWR VPWR _12765_/X sky130_fd_sc_hd__clkbuf_2
X_14504_ _11669_/X _14504_/D VGND VGND VPWR VPWR _14504_/Q sky130_fd_sc_hd__dfxtp_1
X_11716_ _11716_/A VGND VGND VPWR VPWR _11721_/A sky130_fd_sc_hd__clkbuf_2
X_15484_ _15510_/CLK _15484_/D VGND VGND VPWR VPWR wdata[10] sky130_fd_sc_hd__dfxtp_4
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12692_/X _12146_/X _12472_/X _12695_/X VGND VGND VPWR VPWR _12696_/Y sky130_fd_sc_hd__o22ai_1
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14435_ _11905_/X _14435_/D VGND VGND VPWR VPWR _14435_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _11647_/A VGND VGND VPWR VPWR _11647_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14366_ _15662_/CLK pc[27] VGND VGND VPWR VPWR _14366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11578_ _11578_/A VGND VGND VPWR VPWR _11578_/X sky130_fd_sc_hd__buf_1
XFILLER_116_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13317_ _13316_/X _13321_/X _13393_/S VGND VGND VPWR VPWR _13317_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10529_ _10531_/A VGND VGND VPWR VPWR _10529_/X sky130_fd_sc_hd__clkbuf_1
X_14297_ _15604_/CLK _15464_/Q VGND VGND VPWR VPWR _14297_/Q sky130_fd_sc_hd__dfxtp_1
X_13248_ _13303_/X _13302_/X _13393_/S VGND VGND VPWR VPWR _13248_/X sky130_fd_sc_hd__mux2_1
X_13179_ _13178_/X _13220_/X _13393_/S VGND VGND VPWR VPWR _13179_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07740_ _15600_/Q VGND VGND VPWR VPWR _07740_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07671_ _13126_/X VGND VGND VPWR VPWR _07671_/X sky130_fd_sc_hd__buf_1
XFILLER_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09410_ _09410_/A VGND VGND VPWR VPWR _09410_/X sky130_fd_sc_hd__buf_1
XFILLER_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09341_ _15095_/Q _09335_/X _09206_/X _09336_/X VGND VGND VPWR VPWR _15095_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09272_ _15112_/Q _09262_/X _09271_/X _09264_/X VGND VGND VPWR VPWR _15112_/D sky130_fd_sc_hd__a22o_1
X_08223_ _14300_/Q _08223_/B VGND VGND VPWR VPWR _08660_/A sky130_fd_sc_hd__or2_1
X_08154_ _08184_/A VGND VGND VPWR VPWR _08174_/A sky130_fd_sc_hd__buf_2
XFILLER_147_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07105_ _15667_/Q VGND VGND VPWR VPWR _07383_/A sky130_fd_sc_hd__buf_1
XFILLER_107_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08085_ _15398_/Q _08077_/X _08084_/X _08080_/X VGND VGND VPWR VPWR _15398_/D sky130_fd_sc_hd__a22o_1
XFILLER_146_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08987_ _08989_/A VGND VGND VPWR VPWR _08987_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07938_ _11850_/A VGND VGND VPWR VPWR _08191_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_87_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07869_ _07869_/A VGND VGND VPWR VPWR _07869_/X sky130_fd_sc_hd__buf_1
XFILLER_83_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09608_ _15028_/Q _09593_/X _09607_/X _09597_/X VGND VGND VPWR VPWR _15028_/D sky130_fd_sc_hd__a22o_1
X_10880_ _14711_/Q _10874_/X _10728_/X _10875_/X VGND VGND VPWR VPWR _14711_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09539_ _10308_/A VGND VGND VPWR VPWR _09539_/X sky130_fd_sc_hd__buf_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12550_ _15472_/Q VGND VGND VPWR VPWR _12550_/Y sky130_fd_sc_hd__inv_2
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11501_ _11513_/A VGND VGND VPWR VPWR _11501_/X sky130_fd_sc_hd__buf_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _13171_/X _12451_/X _12389_/X _12459_/X _12480_/X VGND VGND VPWR VPWR _12481_/X
+ sky130_fd_sc_hd__o221a_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ _14954_/Q _15050_/Q _15018_/Q _15082_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14220_/X sky130_fd_sc_hd__mux4_2
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11432_ _11446_/A VGND VGND VPWR VPWR _11450_/A sky130_fd_sc_hd__inv_2
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14151_ _14147_/X _14148_/X _14149_/X _14150_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14151_/X sky130_fd_sc_hd__mux4_1
X_11363_ _11393_/A VGND VGND VPWR VPWR _11384_/A sky130_fd_sc_hd__buf_2
XFILLER_138_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13102_ _15648_/Q data_address[13] _15667_/Q VGND VGND VPWR VPWR _13102_/X sky130_fd_sc_hd__mux2_1
X_10314_ _10314_/A VGND VGND VPWR VPWR _10314_/X sky130_fd_sc_hd__clkbuf_2
X_14082_ _15223_/Q _14551_/Q _14999_/Q _15415_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14082_/X sky130_fd_sc_hd__mux4_1
X_11294_ _11303_/A VGND VGND VPWR VPWR _11294_/X sky130_fd_sc_hd__buf_1
XFILLER_98_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13033_ wdata[6] rdata[6] _13058_/S VGND VGND VPWR VPWR _14310_/D sky130_fd_sc_hd__mux2_1
X_10245_ _14865_/Q _10237_/X _10008_/X _10238_/X VGND VGND VPWR VPWR _14865_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10176_ _10180_/A VGND VGND VPWR VPWR _10176_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14984_ _09792_/X _14984_/D VGND VGND VPWR VPWR _14984_/Q sky130_fd_sc_hd__dfxtp_1
X_13935_ _15110_/Q _15334_/Q _15302_/Q _15270_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13935_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13866_ _13862_/X _13863_/X _13864_/X _13865_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13866_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15605_ _15668_/CLK _15605_/D VGND VGND VPWR VPWR pc[0] sky130_fd_sc_hd__dfxtp_1
X_12817_ _13418_/S _12817_/B VGND VGND VPWR VPWR _12926_/B sky130_fd_sc_hd__nor2_2
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13797_ _14644_/Q _14612_/Q _14580_/Q _15380_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13797_/X sky130_fd_sc_hd__mux4_2
XFILLER_90_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15536_ _15578_/CLK _15536_/D VGND VGND VPWR VPWR _15536_/Q sky130_fd_sc_hd__dfxtp_1
X_12748_ _12746_/X _12201_/A _12747_/Y _12277_/A VGND VGND VPWR VPWR _12749_/B sky130_fd_sc_hd__a31o_1
XFILLER_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15467_ _15521_/CLK _15467_/D VGND VGND VPWR VPWR _15467_/Q sky130_fd_sc_hd__dfxtp_1
X_12679_ _12662_/A _12676_/X _12502_/X VGND VGND VPWR VPWR _12679_/Y sky130_fd_sc_hd__o21ai_1
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14418_ _11969_/X _14418_/D VGND VGND VPWR VPWR _14418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15398_ _08082_/X _15398_/D VGND VGND VPWR VPWR _15398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14349_ _15647_/CLK pc[10] VGND VGND VPWR VPWR _14349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater3 _07310_/Y VGND VGND VPWR VPWR _13581_/A1 sky130_fd_sc_hd__buf_8
XFILLER_98_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08910_ _15206_/Q _08904_/X _08909_/X _08906_/X VGND VGND VPWR VPWR _15206_/D sky130_fd_sc_hd__a22o_1
X_09890_ _14957_/Q _09887_/X _09643_/X _09889_/X VGND VGND VPWR VPWR _14957_/D sky130_fd_sc_hd__a22o_1
X_08841_ _08866_/A VGND VGND VPWR VPWR _08841_/X sky130_fd_sc_hd__buf_1
XFILLER_112_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08772_ _08897_/A VGND VGND VPWR VPWR _08858_/A sky130_fd_sc_hd__buf_2
XFILLER_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07723_ _13142_/X VGND VGND VPWR VPWR _07723_/X sky130_fd_sc_hd__buf_1
XFILLER_65_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07654_ _07675_/A VGND VGND VPWR VPWR _07655_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07585_ _07585_/A _13077_/X VGND VGND VPWR VPWR _15492_/D sky130_fd_sc_hd__and2_1
XFILLER_22_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09324_ _09342_/A VGND VGND VPWR VPWR _09331_/A sky130_fd_sc_hd__buf_1
X_09255_ _09255_/A VGND VGND VPWR VPWR _09255_/X sky130_fd_sc_hd__buf_1
X_08206_ _15367_/Q _08204_/X _08079_/X _08205_/X VGND VGND VPWR VPWR _15367_/D sky130_fd_sc_hd__a22o_1
X_09186_ _15132_/Q _09183_/X _09184_/X _09185_/X VGND VGND VPWR VPWR _15132_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08137_ _08139_/A VGND VGND VPWR VPWR _08137_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08068_ _14310_/Q VGND VGND VPWR VPWR _08069_/A sky130_fd_sc_hd__buf_1
XFILLER_135_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10030_ _10399_/A VGND VGND VPWR VPWR _10030_/X sky130_fd_sc_hd__buf_1
XFILLER_49_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11981_ _11981_/A VGND VGND VPWR VPWR _11981_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13720_ _14972_/Q _15068_/Q _15036_/Q _15100_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13720_/X sky130_fd_sc_hd__mux4_2
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10932_ _11140_/A VGND VGND VPWR VPWR _10999_/A sky130_fd_sc_hd__buf_2
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13651_ _13650_/X _13059_/X _14337_/Q VGND VGND VPWR VPWR _13651_/X sky130_fd_sc_hd__mux2_1
X_10863_ _10869_/A VGND VGND VPWR VPWR _10863_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12602_ _15551_/Q VGND VGND VPWR VPWR _12602_/X sky130_fd_sc_hd__buf_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ _13581_/X _14321_/D _15506_/Q VGND VGND VPWR VPWR _13582_/X sky130_fd_sc_hd__mux2_1
X_10794_ _11537_/A VGND VGND VPWR VPWR _10794_/X sky130_fd_sc_hd__buf_1
XFILLER_9_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15321_ _08404_/X _15321_/D VGND VGND VPWR VPWR _15321_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12533_ _12505_/X _12532_/X _12505_/X _12532_/X VGND VGND VPWR VPWR _12534_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15252_ _08720_/X _15252_/D VGND VGND VPWR VPWR _15252_/Q sky130_fd_sc_hd__dfxtp_1
X_12464_ _15590_/Q VGND VGND VPWR VPWR _12473_/A sky130_fd_sc_hd__inv_2
X_14203_ _14667_/Q _15243_/Q _14731_/Q _14699_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14203_/X sky130_fd_sc_hd__mux4_2
X_11415_ _11415_/A VGND VGND VPWR VPWR _11415_/X sky130_fd_sc_hd__buf_1
XFILLER_126_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15183_ _08996_/X _15183_/D VGND VGND VPWR VPWR _15183_/Q sky130_fd_sc_hd__dfxtp_1
X_12395_ _12395_/A _12395_/B VGND VGND VPWR VPWR _12395_/Y sky130_fd_sc_hd__nand2_2
XFILLER_137_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14134_ _15186_/Q _15154_/Q _14770_/Q _14802_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14134_/X sky130_fd_sc_hd__mux4_1
X_11346_ _11439_/A VGND VGND VPWR VPWR _11407_/A sky130_fd_sc_hd__buf_1
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14065_ _15129_/Q _15353_/Q _15321_/Q _15289_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14065_/X sky130_fd_sc_hd__mux4_1
X_11277_ _14607_/Q _11273_/X _11152_/X _11274_/X VGND VGND VPWR VPWR _14607_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13016_ _14360_/Q VGND VGND VPWR VPWR _13016_/Y sky130_fd_sc_hd__inv_2
X_10228_ _10258_/A VGND VGND VPWR VPWR _10248_/A sky130_fd_sc_hd__buf_2
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10159_ _14890_/Q _10157_/X _10038_/X _10158_/X VGND VGND VPWR VPWR _14890_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14967_ _09852_/X _14967_/D VGND VGND VPWR VPWR _14967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13918_ _14504_/Q _14472_/Q _14440_/Q _14408_/Q _13918_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13918_/X sky130_fd_sc_hd__mux4_2
X_14898_ _10130_/X _14898_/D VGND VGND VPWR VPWR _14898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13849_ _14831_/Q _14863_/Q _14895_/Q _14927_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13849_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07370_ _07377_/A _07370_/B VGND VGND VPWR VPWR _15596_/D sky130_fd_sc_hd__nor2_1
X_15519_ _15521_/CLK _15519_/D VGND VGND VPWR VPWR _15519_/Q sky130_fd_sc_hd__dfxtp_1
X_09040_ _09052_/A VGND VGND VPWR VPWR _09041_/A sky130_fd_sc_hd__buf_1
XFILLER_129_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09942_ _10023_/A VGND VGND VPWR VPWR _09972_/A sky130_fd_sc_hd__buf_2
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09873_ _14962_/Q _09868_/X _09617_/X _09869_/X VGND VGND VPWR VPWR _14962_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08824_ _08829_/A VGND VGND VPWR VPWR _08824_/X sky130_fd_sc_hd__clkbuf_1
X_08755_ _15242_/Q _08753_/X _08505_/X _08754_/X VGND VGND VPWR VPWR _15242_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07706_ _07706_/A VGND VGND VPWR VPWR _07706_/X sky130_fd_sc_hd__buf_1
XFILLER_72_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08686_ _08746_/A VGND VGND VPWR VPWR _08705_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07637_ _07641_/A _07637_/B VGND VGND VPWR VPWR _15463_/D sky130_fd_sc_hd__or2_1
XFILLER_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07568_ _07568_/A _13089_/X VGND VGND VPWR VPWR _15504_/D sky130_fd_sc_hd__and2_1
XFILLER_139_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09307_ _09307_/A VGND VGND VPWR VPWR _09318_/A sky130_fd_sc_hd__buf_1
XFILLER_110_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07499_ _14385_/Q VGND VGND VPWR VPWR _12563_/C sky130_fd_sc_hd__inv_2
X_09238_ _15120_/Q _09235_/X _09236_/X _09237_/X VGND VGND VPWR VPWR _15120_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09169_ _09195_/A VGND VGND VPWR VPWR _09169_/X sky130_fd_sc_hd__buf_1
XFILLER_79_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11200_ _11200_/A VGND VGND VPWR VPWR _11200_/X sky130_fd_sc_hd__clkbuf_1
X_12180_ _15572_/Q VGND VGND VPWR VPWR _12755_/A sky130_fd_sc_hd__inv_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11131_ _14644_/Q _11120_/X _11130_/X _11123_/X VGND VGND VPWR VPWR _14644_/D sky130_fd_sc_hd__a22o_1
XFILLER_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11062_ _11317_/A _11062_/B VGND VGND VPWR VPWR _11078_/A sky130_fd_sc_hd__or2_2
XFILLER_103_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10013_ _10013_/A VGND VGND VPWR VPWR _10013_/X sky130_fd_sc_hd__buf_1
XFILLER_0_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14821_ _10427_/X _14821_/D VGND VGND VPWR VPWR _14821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14752_ _10675_/X _14752_/D VGND VGND VPWR VPWR _14752_/Q sky130_fd_sc_hd__dfxtp_1
X_11964_ _11964_/A VGND VGND VPWR VPWR _11971_/A sky130_fd_sc_hd__buf_1
X_13703_ _14685_/Q _15261_/Q _14749_/Q _14717_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13703_/X sky130_fd_sc_hd__mux4_2
X_10915_ _10915_/A VGND VGND VPWR VPWR _10937_/A sky130_fd_sc_hd__buf_1
X_14683_ _10980_/X _14683_/D VGND VGND VPWR VPWR _14683_/Q sky130_fd_sc_hd__dfxtp_1
X_11895_ _11895_/A VGND VGND VPWR VPWR _11895_/X sky130_fd_sc_hd__buf_1
XFILLER_60_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13634_ _13633_/X _14308_/D _15506_/Q VGND VGND VPWR VPWR _13634_/X sky130_fd_sc_hd__mux2_1
X_10846_ _14721_/Q _10840_/X _10672_/X _10843_/X VGND VGND VPWR VPWR _14721_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13565_ _13564_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13565_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10777_ _14734_/Q _10764_/X _10776_/X _10767_/X VGND VGND VPWR VPWR _14734_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15304_ _08514_/X _15304_/D VGND VGND VPWR VPWR _15304_/Q sky130_fd_sc_hd__dfxtp_1
X_12516_ _15560_/Q VGND VGND VPWR VPWR _12522_/A sky130_fd_sc_hd__inv_2
XFILLER_9_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13496_ _13495_/X _13068_/X _14336_/Q VGND VGND VPWR VPWR _13496_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15235_ _08775_/X _15235_/D VGND VGND VPWR VPWR _15235_/Q sky130_fd_sc_hd__dfxtp_1
X_12447_ _12447_/A VGND VGND VPWR VPWR _12447_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15166_ _09060_/X _15166_/D VGND VGND VPWR VPWR _15166_/Q sky130_fd_sc_hd__dfxtp_1
X_12378_ _15555_/Q VGND VGND VPWR VPWR _12379_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_141_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14117_ _14644_/Q _14612_/Q _14580_/Q _15380_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14117_/X sky130_fd_sc_hd__mux4_2
X_11329_ _11329_/A VGND VGND VPWR VPWR _11329_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15097_ _09334_/X _15097_/D VGND VGND VPWR VPWR _15097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14048_ _14523_/Q _14491_/Q _14459_/Q _14427_/Q _14395_/Q _14060_/S1 VGND VGND VPWR
+ VPWR _14048_/X sky130_fd_sc_hd__mux4_2
XFILLER_122_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08540_ _09287_/A VGND VGND VPWR VPWR _08540_/X sky130_fd_sc_hd__buf_1
XFILLER_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08471_ _10770_/A VGND VGND VPWR VPWR _09240_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07422_ _07424_/A _13595_/X VGND VGND VPWR VPWR _15575_/D sky130_fd_sc_hd__and2_1
XFILLER_62_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07353_ _07353_/A _07353_/B VGND VGND VPWR VPWR _15598_/D sky130_fd_sc_hd__nor2_1
X_07284_ _07286_/A _07284_/B VGND VGND VPWR VPWR _15612_/D sky130_fd_sc_hd__nor2_1
XFILLER_148_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09023_ _09023_/A VGND VGND VPWR VPWR _09030_/A sky130_fd_sc_hd__buf_1
XFILLER_105_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09925_ _10838_/A _10181_/B VGND VGND VPWR VPWR _09941_/A sky130_fd_sc_hd__or2_2
XFILLER_132_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09856_ _09877_/A VGND VGND VPWR VPWR _09856_/X sky130_fd_sc_hd__buf_1
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08807_ _08807_/A VGND VGND VPWR VPWR _08816_/A sky130_fd_sc_hd__buf_1
XFILLER_46_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09787_ _09797_/A VGND VGND VPWR VPWR _09787_/X sky130_fd_sc_hd__buf_1
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08738_ _08740_/A VGND VGND VPWR VPWR _08738_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_105 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_116 rdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 rdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 rdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_149 rdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08669_ _08669_/A VGND VGND VPWR VPWR _08669_/X sky130_fd_sc_hd__buf_1
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10700_ _10706_/A VGND VGND VPWR VPWR _10700_/X sky130_fd_sc_hd__clkbuf_1
X_11680_ _11680_/A VGND VGND VPWR VPWR _11685_/A sky130_fd_sc_hd__buf_1
XFILLER_42_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10631_ _10640_/A VGND VGND VPWR VPWR _10636_/A sky130_fd_sc_hd__buf_1
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13350_ _13352_/X _13351_/X _13408_/S VGND VGND VPWR VPWR _13350_/X sky130_fd_sc_hd__mux2_1
X_10562_ _10562_/A VGND VGND VPWR VPWR _10626_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12301_ _12301_/A VGND VGND VPWR VPWR _12437_/A sky130_fd_sc_hd__buf_1
XFILLER_127_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13281_ _13282_/X _13314_/X _13408_/S VGND VGND VPWR VPWR _13281_/X sky130_fd_sc_hd__mux2_1
X_10493_ _10555_/A VGND VGND VPWR VPWR _10512_/A sky130_fd_sc_hd__buf_4
XFILLER_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15020_ _09647_/X _15020_/D VGND VGND VPWR VPWR _15020_/Q sky130_fd_sc_hd__dfxtp_1
X_12232_ _12216_/Y _12863_/A _12228_/Y _12231_/X VGND VGND VPWR VPWR _12800_/A sky130_fd_sc_hd__a31o_1
XFILLER_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12163_ _15541_/Q VGND VGND VPWR VPWR _12720_/A sky130_fd_sc_hd__inv_2
X_11114_ _11128_/A VGND VGND VPWR VPWR _11125_/A sky130_fd_sc_hd__buf_1
XFILLER_123_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12094_ _12094_/A VGND VGND VPWR VPWR _12094_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11045_ _11045_/A VGND VGND VPWR VPWR _11045_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14804_ _10490_/X _14804_/D VGND VGND VPWR VPWR _14804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12996_ _14340_/Q VGND VGND VPWR VPWR _12996_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14735_ _10769_/X _14735_/D VGND VGND VPWR VPWR _14735_/Q sky130_fd_sc_hd__dfxtp_1
X_11947_ _11947_/A VGND VGND VPWR VPWR _11947_/X sky130_fd_sc_hd__buf_1
XFILLER_18_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14666_ _11036_/X _14666_/D VGND VGND VPWR VPWR _14666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11878_ _14445_/Q _11875_/X _08048_/A _11877_/X VGND VGND VPWR VPWR _14445_/D sky130_fd_sc_hd__a22o_1
XFILLER_33_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13617_ _13616_/X _07336_/Y _13641_/S VGND VGND VPWR VPWR _13617_/X sky130_fd_sc_hd__mux2_1
X_10829_ _14724_/Q _10663_/A _10828_/X _10668_/A VGND VGND VPWR VPWR _14724_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14597_ _11308_/X _14597_/D VGND VGND VPWR VPWR _14597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13548_ _14036_/X _14041_/X _14387_/Q VGND VGND VPWR VPWR _13548_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13479_ _13826_/X _13831_/X _13521_/S VGND VGND VPWR VPWR _13479_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15218_ _08855_/X _15218_/D VGND VGND VPWR VPWR _15218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15149_ _09114_/X _15149_/D VGND VGND VPWR VPWR _15149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07971_ _07971_/A VGND VGND VPWR VPWR _07971_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09710_ _15008_/Q _09702_/X _09539_/X _09705_/X VGND VGND VPWR VPWR _15008_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09641_ _09675_/A VGND VGND VPWR VPWR _09641_/X sky130_fd_sc_hd__buf_1
XFILLER_110_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09572_ _09582_/A VGND VGND VPWR VPWR _09572_/X sky130_fd_sc_hd__clkbuf_1
X_08523_ _09275_/A VGND VGND VPWR VPWR _08523_/X sky130_fd_sc_hd__buf_1
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08454_ _09228_/A VGND VGND VPWR VPWR _08454_/X sky130_fd_sc_hd__buf_1
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07405_ _07406_/A _13551_/X VGND VGND VPWR VPWR _15586_/D sky130_fd_sc_hd__and2_1
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08385_ _15325_/Q _08366_/X _08384_/X _08372_/X VGND VGND VPWR VPWR _15325_/D sky130_fd_sc_hd__a22o_1
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07336_ _07337_/B VGND VGND VPWR VPWR _07336_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07267_ _07269_/A _07267_/B VGND VGND VPWR VPWR _15624_/D sky130_fd_sc_hd__nor2_1
X_09006_ _09025_/A VGND VGND VPWR VPWR _09006_/X sky130_fd_sc_hd__buf_1
XFILLER_124_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07198_ _07209_/A VGND VGND VPWR VPWR _07198_/X sky130_fd_sc_hd__buf_1
XFILLER_145_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09908_ _09908_/A VGND VGND VPWR VPWR _09908_/X sky130_fd_sc_hd__buf_1
X_09839_ _14972_/Q _09837_/X _09564_/X _09838_/X VGND VGND VPWR VPWR _14972_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12850_ _12850_/A _12883_/A VGND VGND VPWR VPWR _12851_/A sky130_fd_sc_hd__or2_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11801_ _11811_/A VGND VGND VPWR VPWR _11814_/A sky130_fd_sc_hd__inv_2
X_12781_ _12778_/X _12204_/X _12753_/X _12780_/X VGND VGND VPWR VPWR _12781_/Y sky130_fd_sc_hd__o22ai_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14520_ _11615_/X _14520_/D VGND VGND VPWR VPWR _14520_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11732_ _11763_/A VGND VGND VPWR VPWR _11752_/A sky130_fd_sc_hd__clkbuf_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14451_ _11855_/X _14451_/D VGND VGND VPWR VPWR _14451_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11663_ _11669_/A VGND VGND VPWR VPWR _11663_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13402_ _13404_/X _13403_/X _13415_/S VGND VGND VPWR VPWR _13402_/X sky130_fd_sc_hd__mux2_1
X_10614_ _14769_/Q _10607_/X _10375_/X _10608_/X VGND VGND VPWR VPWR _14769_/D sky130_fd_sc_hd__a22o_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14382_ _14392_/CLK instruction[11] VGND VGND VPWR VPWR _14382_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ _11613_/A VGND VGND VPWR VPWR _11594_/X sky130_fd_sc_hd__buf_1
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13333_ _13373_/X _13371_/X _13415_/S VGND VGND VPWR VPWR _13333_/X sky130_fd_sc_hd__mux2_1
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10545_ _10547_/A VGND VGND VPWR VPWR _10545_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13264_ _13265_/X _13277_/X _15562_/Q VGND VGND VPWR VPWR _13264_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10476_ _14809_/Q _10474_/X _10340_/X _10475_/X VGND VGND VPWR VPWR _14809_/D sky130_fd_sc_hd__a22o_1
X_15003_ _09729_/X _15003_/D VGND VGND VPWR VPWR _15003_/Q sky130_fd_sc_hd__dfxtp_1
X_12215_ _12230_/A _12230_/B VGND VGND VPWR VPWR _12215_/Y sky130_fd_sc_hd__nor2_2
XFILLER_123_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13195_ _13194_/X _13280_/X _15565_/Q VGND VGND VPWR VPWR _13195_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12146_ _15576_/Q VGND VGND VPWR VPWR _12146_/X sky130_fd_sc_hd__buf_1
XFILLER_96_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12077_ _12577_/A _12075_/B _12586_/A VGND VGND VPWR VPWR _12598_/A sky130_fd_sc_hd__a21oi_2
XFILLER_110_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11028_ _14669_/Q _11025_/X _10782_/X _11027_/X VGND VGND VPWR VPWR _14669_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12979_ _12979_/A _12979_/B VGND VGND VPWR VPWR _13076_/S sky130_fd_sc_hd__nor2_8
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14718_ _10858_/X _14718_/D VGND VGND VPWR VPWR _14718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14649_ _11106_/X _14649_/D VGND VGND VPWR VPWR _14649_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_16 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_27 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08170_ _15377_/Q _08164_/X _08026_/X _08165_/X VGND VGND VPWR VPWR _15377_/D sky130_fd_sc_hd__a22o_1
XANTENNA_38 data_address[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 data_address[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07121_ _12023_/D VGND VGND VPWR VPWR _12040_/B sky130_fd_sc_hd__buf_1
XFILLER_119_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07954_ _07984_/A VGND VGND VPWR VPWR _07954_/X sky130_fd_sc_hd__buf_1
XFILLER_68_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07885_ _07885_/A VGND VGND VPWR VPWR _07885_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09624_ _09630_/A VGND VGND VPWR VPWR _09624_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09555_ _09603_/A VGND VGND VPWR VPWR _09586_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08506_ _08524_/A VGND VGND VPWR VPWR _08506_/X sky130_fd_sc_hd__buf_1
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09486_ _09505_/A VGND VGND VPWR VPWR _09486_/X sky130_fd_sc_hd__buf_1
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08437_ _08547_/A VGND VGND VPWR VPWR _08474_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08368_ _10683_/A VGND VGND VPWR VPWR _09170_/A sky130_fd_sc_hd__buf_1
X_07319_ _07319_/A VGND VGND VPWR VPWR _07319_/X sky130_fd_sc_hd__buf_1
XFILLER_149_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08299_ _08319_/A VGND VGND VPWR VPWR _08304_/A sky130_fd_sc_hd__buf_2
X_10330_ _14844_/Q _10327_/X _10328_/X _10329_/X VGND VGND VPWR VPWR _14844_/D sky130_fd_sc_hd__a22o_1
XFILLER_125_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10261_ _10261_/A VGND VGND VPWR VPWR _10266_/A sky130_fd_sc_hd__buf_1
XFILLER_152_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12000_ _14409_/Q _11996_/X _08069_/A _11997_/X VGND VGND VPWR VPWR _14409_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10192_ _14880_/Q _10183_/X _09938_/X _10186_/X VGND VGND VPWR VPWR _14880_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13951_ _13947_/X _13948_/X _13949_/X _13950_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13951_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12902_ _12902_/A _12902_/B _12902_/C VGND VGND VPWR VPWR _12902_/X sky130_fd_sc_hd__or3_1
XFILLER_86_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13882_ _15211_/Q _14539_/Q _14987_/Q _15403_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13882_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15621_ _15621_/CLK _15621_/D VGND VGND VPWR VPWR pc[16] sky130_fd_sc_hd__dfxtp_4
X_12833_ _12802_/A _12802_/B _12428_/A _12803_/B VGND VGND VPWR VPWR _12833_/Y sky130_fd_sc_hd__o211ai_4
X_12764_ _12762_/X _12763_/X _12677_/X _13273_/X _12710_/X VGND VGND VPWR VPWR _12764_/X
+ sky130_fd_sc_hd__o32a_1
X_15552_ _15590_/CLK _15552_/D VGND VGND VPWR VPWR _15552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14503_ _11672_/X _14503_/D VGND VGND VPWR VPWR _14503_/Q sky130_fd_sc_hd__dfxtp_1
X_11715_ _14492_/Q _11713_/X _11463_/X _11714_/X VGND VGND VPWR VPWR _14492_/D sky130_fd_sc_hd__a22o_1
X_15483_ _15521_/CLK _15483_/D VGND VGND VPWR VPWR wdata[9] sky130_fd_sc_hd__dfxtp_2
X_12695_ _12703_/A _12703_/B _12475_/X VGND VGND VPWR VPWR _12695_/X sky130_fd_sc_hd__o21a_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11646_ _14511_/Q _11642_/X _11518_/X _11643_/X VGND VGND VPWR VPWR _14511_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14434_ _11909_/X _14434_/D VGND VGND VPWR VPWR _14434_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ _15663_/CLK pc[26] VGND VGND VPWR VPWR _14365_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11577_ _11589_/A VGND VGND VPWR VPWR _11578_/A sky130_fd_sc_hd__buf_1
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13316_ _13415_/X _13412_/X _13408_/S VGND VGND VPWR VPWR _13316_/X sky130_fd_sc_hd__mux2_1
X_10528_ _14794_/Q _10526_/X _10407_/X _10527_/X VGND VGND VPWR VPWR _14794_/D sky130_fd_sc_hd__a22o_1
X_14296_ _15510_/CLK _15463_/Q VGND VGND VPWR VPWR _14296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13247_ _12709_/X _12730_/A _13418_/S VGND VGND VPWR VPWR _13247_/X sky130_fd_sc_hd__mux2_1
X_10459_ _14814_/Q _10453_/X _10320_/X _10456_/X VGND VGND VPWR VPWR _14814_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13178_ _13181_/X _13201_/X _13408_/S VGND VGND VPWR VPWR _13178_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12129_ _12148_/A VGND VGND VPWR VPWR _12130_/A sky130_fd_sc_hd__buf_1
XFILLER_69_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07670_ _07781_/A VGND VGND VPWR VPWR _07670_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09340_ _09340_/A VGND VGND VPWR VPWR _09340_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09271_ _09271_/A VGND VGND VPWR VPWR _09271_/X sky130_fd_sc_hd__buf_1
XFILLER_21_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08222_ _08550_/B VGND VGND VPWR VPWR _09150_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08153_ _08173_/A VGND VGND VPWR VPWR _08153_/X sky130_fd_sc_hd__buf_1
XFILLER_119_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08084_ _08084_/A VGND VGND VPWR VPWR _08084_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08986_ _15187_/Q _08984_/X _08852_/X _08985_/X VGND VGND VPWR VPWR _15187_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07937_ _15425_/Q _07927_/X _07936_/X _07932_/X VGND VGND VPWR VPWR _15425_/D sky130_fd_sc_hd__a22o_1
X_07868_ _07868_/A VGND VGND VPWR VPWR _07868_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09607_ _10363_/A VGND VGND VPWR VPWR _09607_/X sky130_fd_sc_hd__buf_1
X_07799_ _07659_/X _07664_/X _07798_/X VGND VGND VPWR VPWR _07800_/A sky130_fd_sc_hd__o21ai_1
XFILLER_71_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09538_ _10676_/A VGND VGND VPWR VPWR _10308_/A sky130_fd_sc_hd__buf_1
XFILLER_71_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09469_ _09469_/A VGND VGND VPWR VPWR _09474_/A sky130_fd_sc_hd__buf_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11500_ _11505_/A VGND VGND VPWR VPWR _11500_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12480_ _12480_/A _12480_/B _12789_/A VGND VGND VPWR VPWR _12480_/X sky130_fd_sc_hd__or3_2
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11431_ _11431_/A VGND VGND VPWR VPWR _11431_/X sky130_fd_sc_hd__buf_1
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14150_ _14961_/Q _15057_/Q _15025_/Q _15089_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14150_/X sky130_fd_sc_hd__mux4_1
X_11362_ _11362_/A VGND VGND VPWR VPWR _11362_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13101_ _15647_/Q data_address[12] _15667_/Q VGND VGND VPWR VPWR _13101_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10313_ _10339_/A VGND VGND VPWR VPWR _10313_/X sky130_fd_sc_hd__buf_1
XFILLER_125_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14081_ _14077_/X _14078_/X _14079_/X _14080_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14081_/X sky130_fd_sc_hd__mux4_1
X_11293_ _11299_/A VGND VGND VPWR VPWR _11293_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13032_ wdata[5] rdata[5] _13058_/S VGND VGND VPWR VPWR _14309_/D sky130_fd_sc_hd__mux2_4
XFILLER_106_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10244_ _10246_/A VGND VGND VPWR VPWR _10244_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10175_ _10201_/A VGND VGND VPWR VPWR _10180_/A sky130_fd_sc_hd__buf_1
XFILLER_120_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14983_ _09796_/X _14983_/D VGND VGND VPWR VPWR _14983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13934_ _15174_/Q _15142_/Q _14758_/Q _14790_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13934_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13865_ _15117_/Q _15341_/Q _15309_/Q _15277_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13865_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15604_ _15604_/CLK _15604_/D VGND VGND VPWR VPWR _15604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12816_ _15529_/Q VGND VGND VPWR VPWR _12817_/B sky130_fd_sc_hd__clkinv_4
X_13796_ _13792_/X _13793_/X _13794_/X _13795_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13796_/X sky130_fd_sc_hd__mux4_2
XFILLER_15_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15535_ _15566_/CLK _15535_/D VGND VGND VPWR VPWR _15535_/Q sky130_fd_sc_hd__dfxtp_1
X_12747_ _12747_/A VGND VGND VPWR VPWR _12747_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _12662_/X _12676_/X _12677_/X _13393_/X _12496_/X VGND VGND VPWR VPWR _12678_/X
+ sky130_fd_sc_hd__o32a_1
X_15466_ _15509_/CLK _15466_/D VGND VGND VPWR VPWR _15466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14417_ _11971_/X _14417_/D VGND VGND VPWR VPWR _14417_/Q sky130_fd_sc_hd__dfxtp_1
X_11629_ _14516_/Q _11622_/X _11498_/X _11624_/X VGND VGND VPWR VPWR _14516_/D sky130_fd_sc_hd__a22o_1
X_15397_ _08089_/X _15397_/D VGND VGND VPWR VPWR _15397_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14348_ _15646_/CLK pc[9] VGND VGND VPWR VPWR _14348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14279_ _14820_/Q _14852_/Q _14884_/Q _14916_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14279_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater4 _13641_/S VGND VGND VPWR VPWR _13569_/S sky130_fd_sc_hd__buf_8
XFILLER_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08840_ _08879_/A VGND VGND VPWR VPWR _08866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08771_ _15236_/Q _08666_/A _08540_/X _08669_/A VGND VGND VPWR VPWR _15236_/D sky130_fd_sc_hd__a22o_1
X_07722_ _07722_/A VGND VGND VPWR VPWR _07772_/A sky130_fd_sc_hd__inv_2
XFILLER_26_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07653_ _07653_/A VGND VGND VPWR VPWR _07675_/A sky130_fd_sc_hd__buf_1
XFILLER_81_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07584_ _07585_/A _13078_/X VGND VGND VPWR VPWR _15493_/D sky130_fd_sc_hd__and2_1
XFILLER_80_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09323_ _09383_/A VGND VGND VPWR VPWR _09342_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09254_ _09254_/A VGND VGND VPWR VPWR _09254_/X sky130_fd_sc_hd__clkbuf_1
X_08205_ _08205_/A VGND VGND VPWR VPWR _08205_/X sky130_fd_sc_hd__buf_1
XFILLER_21_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09185_ _09197_/A VGND VGND VPWR VPWR _09185_/X sky130_fd_sc_hd__buf_1
XFILLER_147_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08136_ _15388_/Q _08134_/X _07968_/X _08135_/X VGND VGND VPWR VPWR _15388_/D sky130_fd_sc_hd__a22o_1
XFILLER_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08067_ _08067_/A VGND VGND VPWR VPWR _08067_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08969_ _15191_/Q _08963_/X _08834_/X _08964_/X VGND VGND VPWR VPWR _15191_/D sky130_fd_sc_hd__a22o_1
X_11980_ _14415_/Q _11976_/X _08036_/A _11977_/X VGND VGND VPWR VPWR _14415_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10931_ _10931_/A VGND VGND VPWR VPWR _11140_/A sky130_fd_sc_hd__buf_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10862_ _10862_/A VGND VGND VPWR VPWR _10869_/A sky130_fd_sc_hd__buf_1
X_13650_ _13649_/X _14304_/D _15506_/Q VGND VGND VPWR VPWR _13650_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _12599_/X _12577_/X _12600_/X _13301_/X _12319_/X VGND VGND VPWR VPWR _12601_/X
+ sky130_fd_sc_hd__o32a_1
X_13581_ _13580_/X _13581_/A1 _13641_/S VGND VGND VPWR VPWR _13581_/X sky130_fd_sc_hd__mux2_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10793_ _10793_/A VGND VGND VPWR VPWR _11537_/A sky130_fd_sc_hd__clkbuf_2
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15320_ _08411_/X _15320_/D VGND VGND VPWR VPWR _15320_/Q sky130_fd_sc_hd__dfxtp_1
X_12532_ _12951_/C VGND VGND VPWR VPWR _12532_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12463_ _15590_/Q VGND VGND VPWR VPWR _12463_/X sky130_fd_sc_hd__buf_1
X_15251_ _08722_/X _15251_/D VGND VGND VPWR VPWR _15251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11414_ _11414_/A VGND VGND VPWR VPWR _11414_/X sky130_fd_sc_hd__buf_1
X_14202_ _15211_/Q _14539_/Q _14987_/Q _15403_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14202_/X sky130_fd_sc_hd__mux4_1
X_15182_ _08998_/X _15182_/D VGND VGND VPWR VPWR _15182_/Q sky130_fd_sc_hd__dfxtp_1
X_12394_ _12394_/A VGND VGND VPWR VPWR _12432_/A sky130_fd_sc_hd__inv_2
XFILLER_153_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14133_ _14674_/Q _15250_/Q _14738_/Q _14706_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14133_/X sky130_fd_sc_hd__mux4_2
X_11345_ _14588_/Q _11343_/X _11095_/X _11344_/X VGND VGND VPWR VPWR _14588_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14064_ _15193_/Q _15161_/Q _14777_/Q _14809_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14064_/X sky130_fd_sc_hd__mux4_2
XFILLER_4_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11276_ _11278_/A VGND VGND VPWR VPWR _11276_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13015_ _14359_/Q VGND VGND VPWR VPWR _13015_/Y sky130_fd_sc_hd__inv_2
X_10227_ _10247_/A VGND VGND VPWR VPWR _10227_/X sky130_fd_sc_hd__buf_1
XFILLER_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10158_ _10167_/A VGND VGND VPWR VPWR _10158_/X sky130_fd_sc_hd__buf_1
XFILLER_0_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14966_ _09854_/X _14966_/D VGND VGND VPWR VPWR _14966_/Q sky130_fd_sc_hd__dfxtp_1
X_10089_ _10107_/A VGND VGND VPWR VPWR _10089_/X sky130_fd_sc_hd__buf_1
XFILLER_94_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13917_ _14632_/Q _14600_/Q _14568_/Q _15368_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13917_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14897_ _10132_/X _14897_/D VGND VGND VPWR VPWR _14897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13848_ _14511_/Q _14479_/Q _14447_/Q _14415_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13848_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13779_ _14838_/Q _14870_/Q _14902_/Q _14934_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13779_/X sky130_fd_sc_hd__mux4_2
XFILLER_50_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15518_ _15521_/CLK _15518_/D VGND VGND VPWR VPWR _15518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15449_ _15647_/CLK _15449_/D VGND VGND VPWR VPWR data_address[22] sky130_fd_sc_hd__dfxtp_4
XFILLER_129_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09941_ _09941_/A VGND VGND VPWR VPWR _10023_/A sky130_fd_sc_hd__clkbuf_2
X_09872_ _09876_/A VGND VGND VPWR VPWR _09872_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08823_ _15226_/Q _08812_/X _08822_/X _08814_/X VGND VGND VPWR VPWR _15226_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08754_ _08763_/A VGND VGND VPWR VPWR _08754_/X sky130_fd_sc_hd__buf_1
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07705_ _07705_/A VGND VGND VPWR VPWR _07777_/B sky130_fd_sc_hd__inv_2
XFILLER_26_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08685_ _08897_/A VGND VGND VPWR VPWR _08746_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07636_ _15511_/Q VGND VGND VPWR VPWR _07637_/B sky130_fd_sc_hd__buf_1
XFILLER_81_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07567_ _07568_/A _13090_/X VGND VGND VPWR VPWR _15505_/D sky130_fd_sc_hd__and2_1
X_09306_ _15104_/Q _09298_/X _09164_/X _09301_/X VGND VGND VPWR VPWR _15104_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07498_ _07500_/A _07498_/B VGND VGND VPWR VPWR _15522_/D sky130_fd_sc_hd__nor2_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09237_ _09237_/A VGND VGND VPWR VPWR _09237_/X sky130_fd_sc_hd__buf_1
X_09168_ _09248_/A VGND VGND VPWR VPWR _09195_/A sky130_fd_sc_hd__buf_2
XFILLER_107_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08119_ _08129_/A VGND VGND VPWR VPWR _08119_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09099_ _09161_/A VGND VGND VPWR VPWR _09120_/A sky130_fd_sc_hd__buf_2
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11130_ _11498_/A VGND VGND VPWR VPWR _11130_/X sky130_fd_sc_hd__buf_1
XFILLER_134_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11061_ _11061_/A VGND VGND VPWR VPWR _11317_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_89_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10012_ _10379_/A VGND VGND VPWR VPWR _10012_/X sky130_fd_sc_hd__buf_1
XFILLER_88_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14820_ _10430_/X _14820_/D VGND VGND VPWR VPWR _14820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14751_ _10679_/X _14751_/D VGND VGND VPWR VPWR _14751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11963_ _14420_/Q _11956_/X _08011_/A _11958_/X VGND VGND VPWR VPWR _14420_/D sky130_fd_sc_hd__a22o_1
XFILLER_45_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13702_ _15229_/Q _14557_/Q _15005_/Q _15421_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13702_/X sky130_fd_sc_hd__mux4_1
X_10914_ _10936_/A VGND VGND VPWR VPWR _10914_/X sky130_fd_sc_hd__buf_1
XFILLER_17_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14682_ _10982_/X _14682_/D VGND VGND VPWR VPWR _14682_/Q sky130_fd_sc_hd__dfxtp_1
X_11894_ _11898_/A VGND VGND VPWR VPWR _11894_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13633_ _13632_/X _07360_/Y _13641_/S VGND VGND VPWR VPWR _13633_/X sky130_fd_sc_hd__mux2_1
X_10845_ _10847_/A VGND VGND VPWR VPWR _10845_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10776_ _11523_/A VGND VGND VPWR VPWR _10776_/X sky130_fd_sc_hd__buf_1
X_13564_ _14076_/X _14081_/X _13648_/S VGND VGND VPWR VPWR _13564_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15303_ _08519_/X _15303_/D VGND VGND VPWR VPWR _15303_/Q sky130_fd_sc_hd__dfxtp_1
X_12515_ _13167_/X _12493_/X _12497_/X _12504_/Y _12514_/Y VGND VGND VPWR VPWR _12515_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_13495_ _13494_/X rdata[9] _13516_/S VGND VGND VPWR VPWR _13495_/X sky130_fd_sc_hd__mux2_2
XFILLER_9_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12446_ _12902_/A _12446_/B VGND VGND VPWR VPWR _12447_/A sky130_fd_sc_hd__or2_1
X_15234_ _08777_/X _15234_/D VGND VGND VPWR VPWR _15234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12377_ _15587_/Q VGND VGND VPWR VPWR _12379_/A sky130_fd_sc_hd__buf_1
X_15165_ _09062_/X _15165_/D VGND VGND VPWR VPWR _15165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14116_ _14112_/X _14113_/X _14114_/X _14115_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14116_/X sky130_fd_sc_hd__mux4_2
X_11328_ _14592_/Q _11319_/X _11075_/X _11322_/X VGND VGND VPWR VPWR _14592_/D sky130_fd_sc_hd__a22o_1
X_15096_ _09338_/X _15096_/D VGND VGND VPWR VPWR _15096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11259_ _14613_/Q _11254_/X _11126_/X _11256_/X VGND VGND VPWR VPWR _14613_/D sky130_fd_sc_hd__a22o_1
X_14047_ _14651_/Q _14619_/Q _14587_/Q _15387_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14047_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14949_ _09913_/X _14949_/D VGND VGND VPWR VPWR _14949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08470_ _14316_/Q VGND VGND VPWR VPWR _10770_/A sky130_fd_sc_hd__buf_1
XFILLER_35_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07421_ _07429_/A VGND VGND VPWR VPWR _07424_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07352_ _07353_/B VGND VGND VPWR VPWR _07352_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07283_ _07283_/A VGND VGND VPWR VPWR _07286_/A sky130_fd_sc_hd__buf_1
X_09022_ _15176_/Q _09016_/X _08901_/X _09017_/X VGND VGND VPWR VPWR _15176_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09924_ _10294_/B VGND VGND VPWR VPWR _10181_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_131_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09855_ _09886_/A VGND VGND VPWR VPWR _09877_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08806_ _15230_/Q _08798_/X _08805_/X _08802_/X VGND VGND VPWR VPWR _15230_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09786_ _09792_/A VGND VGND VPWR VPWR _09786_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08737_ _15247_/Q _08732_/X _08472_/X _08733_/X VGND VGND VPWR VPWR _15247_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_106 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_117 rdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 rdata[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 rdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08668_ _08680_/A VGND VGND VPWR VPWR _08669_/A sky130_fd_sc_hd__buf_1
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07619_ _07626_/A _07619_/B VGND VGND VPWR VPWR _15473_/D sky130_fd_sc_hd__nor2_1
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08599_ _08618_/A VGND VGND VPWR VPWR _08599_/X sky130_fd_sc_hd__buf_1
XFILLER_81_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10630_ _14765_/Q _10627_/X _10394_/X _10629_/X VGND VGND VPWR VPWR _14765_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10561_ _10561_/A VGND VGND VPWR VPWR _10561_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12300_ _12300_/A VGND VGND VPWR VPWR _12301_/A sky130_fd_sc_hd__buf_1
XFILLER_6_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13280_ _13281_/X _12967_/B _13393_/S VGND VGND VPWR VPWR _13280_/X sky130_fd_sc_hd__mux2_2
X_10492_ _10492_/A VGND VGND VPWR VPWR _10555_/A sky130_fd_sc_hd__buf_1
XFILLER_108_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12231_ _12929_/B _12220_/Y _12230_/Y _12215_/Y VGND VGND VPWR VPWR _12231_/X sky130_fd_sc_hd__a31o_1
XFILLER_108_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12162_ _12162_/A _12689_/A VGND VGND VPWR VPWR _12162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11113_ _14648_/Q _11107_/X _11112_/X _11109_/X VGND VGND VPWR VPWR _14648_/D sky130_fd_sc_hd__a22o_1
XFILLER_150_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12093_ _15581_/Q VGND VGND VPWR VPWR _12627_/A sky130_fd_sc_hd__inv_2
XFILLER_96_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11044_ _14664_/Q _11037_/X _10809_/X _11038_/X VGND VGND VPWR VPWR _14664_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14803_ _10495_/X _14803_/D VGND VGND VPWR VPWR _14803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12995_ _14339_/Q VGND VGND VPWR VPWR _12995_/Y sky130_fd_sc_hd__inv_2
X_14734_ _10774_/X _14734_/D VGND VGND VPWR VPWR _14734_/Q sky130_fd_sc_hd__dfxtp_1
X_11946_ _11946_/A VGND VGND VPWR VPWR _11946_/X sky130_fd_sc_hd__buf_1
XFILLER_17_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14665_ _11041_/X _14665_/D VGND VGND VPWR VPWR _14665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11877_ _11896_/A VGND VGND VPWR VPWR _11877_/X sky130_fd_sc_hd__buf_1
XFILLER_60_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13616_ _14206_/X _14211_/X _13648_/S VGND VGND VPWR VPWR _13616_/X sky130_fd_sc_hd__mux2_2
X_10828_ _11567_/A VGND VGND VPWR VPWR _10828_/X sky130_fd_sc_hd__buf_1
X_14596_ _11312_/X _14596_/D VGND VGND VPWR VPWR _14596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13547_ _13546_/X _13085_/X _14337_/Q VGND VGND VPWR VPWR _13547_/X sky130_fd_sc_hd__mux2_1
X_10759_ _10769_/A VGND VGND VPWR VPWR _10759_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13478_ _13477_/X _13074_/X _14336_/Q VGND VGND VPWR VPWR _13478_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15217_ _08860_/X _15217_/D VGND VGND VPWR VPWR _15217_/Q sky130_fd_sc_hd__dfxtp_1
X_12429_ _12412_/X _12407_/Y _12410_/A VGND VGND VPWR VPWR _12429_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15148_ _09121_/X _15148_/D VGND VGND VPWR VPWR _15148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07970_ _15420_/Q _07966_/X _07968_/X _07969_/X VGND VGND VPWR VPWR _15420_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15079_ _09394_/X _15079_/D VGND VGND VPWR VPWR _15079_/Q sky130_fd_sc_hd__dfxtp_1
X_09640_ _09640_/A VGND VGND VPWR VPWR _09675_/A sky130_fd_sc_hd__buf_1
XFILLER_28_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09571_ _09586_/A VGND VGND VPWR VPWR _09582_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_47_clk _14315_/CLK VGND VGND VPWR VPWR _15647_/CLK sky130_fd_sc_hd__clkbuf_16
X_08522_ _10813_/A VGND VGND VPWR VPWR _09275_/A sky130_fd_sc_hd__buf_1
XFILLER_24_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ _10755_/A VGND VGND VPWR VPWR _09228_/A sky130_fd_sc_hd__buf_1
XFILLER_51_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07404_ _07406_/A _13547_/X VGND VGND VPWR VPWR _15587_/D sky130_fd_sc_hd__and2_1
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08384_ _09180_/A VGND VGND VPWR VPWR _08384_/X sky130_fd_sc_hd__buf_1
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07335_ _07493_/B _07319_/X _07494_/B _07324_/X VGND VGND VPWR VPWR _07337_/B sky130_fd_sc_hd__o22a_1
X_07266_ _07270_/A VGND VGND VPWR VPWR _07269_/A sky130_fd_sc_hd__buf_1
XFILLER_136_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09005_ _09005_/A VGND VGND VPWR VPWR _09025_/A sky130_fd_sc_hd__clkbuf_2
X_07197_ _07197_/A VGND VGND VPWR VPWR _07197_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09907_ _09907_/A VGND VGND VPWR VPWR _09907_/X sky130_fd_sc_hd__buf_1
XFILLER_116_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09838_ _09847_/A VGND VGND VPWR VPWR _09838_/X sky130_fd_sc_hd__buf_1
XFILLER_59_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09769_ _14992_/Q _09767_/X _09627_/X _09768_/X VGND VGND VPWR VPWR _14992_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_38_clk clkbuf_opt_6_clk/X VGND VGND VPWR VPWR _15521_/CLK sky130_fd_sc_hd__clkbuf_16
X_11800_ _11800_/A VGND VGND VPWR VPWR _11800_/X sky130_fd_sc_hd__buf_1
XFILLER_132_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12780_ _12785_/A _12785_/B _12727_/X VGND VGND VPWR VPWR _12780_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11731_ _11731_/A VGND VGND VPWR VPWR _11731_/X sky130_fd_sc_hd__clkbuf_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14450_ _11859_/X _14450_/D VGND VGND VPWR VPWR _14450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11662_ _11680_/A VGND VGND VPWR VPWR _11669_/A sky130_fd_sc_hd__buf_1
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13405_/X _13402_/X _13408_/S VGND VGND VPWR VPWR _13401_/X sky130_fd_sc_hd__mux2_1
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ _10615_/A VGND VGND VPWR VPWR _10613_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14381_ _14381_/CLK instruction[10] VGND VGND VPWR VPWR _14381_/Q sky130_fd_sc_hd__dfxtp_2
X_11593_ _11653_/A VGND VGND VPWR VPWR _11613_/A sky130_fd_sc_hd__buf_2
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13332_ _13370_/X _13367_/X _13415_/S VGND VGND VPWR VPWR _13332_/X sky130_fd_sc_hd__mux2_1
X_10544_ _14788_/Q _10440_/A _10431_/X _10443_/A VGND VGND VPWR VPWR _14788_/D sky130_fd_sc_hd__a22o_1
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13263_ _13264_/X _13287_/X _15563_/Q VGND VGND VPWR VPWR _13263_/X sky130_fd_sc_hd__mux2_1
X_10475_ _10475_/A VGND VGND VPWR VPWR _10475_/X sky130_fd_sc_hd__buf_1
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15002_ _09731_/X _15002_/D VGND VGND VPWR VPWR _15002_/Q sky130_fd_sc_hd__dfxtp_1
X_12214_ _12867_/A _12092_/X _12213_/Y _12094_/X VGND VGND VPWR VPWR _12230_/B sky130_fd_sc_hd__o22a_2
X_13194_ _13193_/X _13235_/X _13393_/S VGND VGND VPWR VPWR _13194_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12145_ _15544_/Q VGND VGND VPWR VPWR _12692_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12076_ _12076_/A VGND VGND VPWR VPWR _12586_/A sky130_fd_sc_hd__inv_2
XFILLER_104_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11027_ _11047_/A VGND VGND VPWR VPWR _11027_/X sky130_fd_sc_hd__buf_1
XFILLER_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clk _14397_/CLK VGND VGND VPWR VPWR _15652_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12978_ _12984_/A _12978_/B VGND VGND VPWR VPWR _13419_/S sky130_fd_sc_hd__nor2_1
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14717_ _10860_/X _14717_/D VGND VGND VPWR VPWR _14717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11929_ _14431_/Q _11925_/X _07951_/A _11928_/X VGND VGND VPWR VPWR _14431_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14648_ _11111_/X _14648_/D VGND VGND VPWR VPWR _14648_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_17 data_address[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_28 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 data_address[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14579_ _11373_/X _14579_/D VGND VGND VPWR VPWR _14579_/Q sky130_fd_sc_hd__dfxtp_1
X_07120_ _15510_/Q _15509_/Q _15508_/Q _15507_/Q VGND VGND VPWR VPWR _12023_/D sky130_fd_sc_hd__or4bb_4
XFILLER_9_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07953_ _08049_/A VGND VGND VPWR VPWR _07984_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07884_ _07884_/A _07884_/B VGND VGND VPWR VPWR _07885_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09623_ _15025_/Q _09610_/X _09622_/X _09613_/X VGND VGND VPWR VPWR _15025_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09554_ _15038_/Q _09544_/X _09553_/X _09549_/X VGND VGND VPWR VPWR _15038_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08505_ _09263_/A VGND VGND VPWR VPWR _08505_/X sky130_fd_sc_hd__buf_1
XFILLER_36_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09485_ _09485_/A VGND VGND VPWR VPWR _09505_/A sky130_fd_sc_hd__buf_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08436_ _08583_/A VGND VGND VPWR VPWR _08547_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08367_ _14332_/Q VGND VGND VPWR VPWR _10683_/A sky130_fd_sc_hd__buf_1
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07318_ _07338_/A VGND VGND VPWR VPWR _07319_/A sky130_fd_sc_hd__buf_1
XFILLER_20_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08298_ _08379_/A VGND VGND VPWR VPWR _08319_/A sky130_fd_sc_hd__buf_1
XFILLER_137_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07249_ _07257_/A VGND VGND VPWR VPWR _07252_/A sky130_fd_sc_hd__clkbuf_2
X_10260_ _14861_/Q _10257_/X _10025_/X _10259_/X VGND VGND VPWR VPWR _14861_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10191_ _10193_/A VGND VGND VPWR VPWR _10191_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13950_ _14949_/Q _15045_/Q _15013_/Q _15077_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13950_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12901_ _12414_/X _12412_/X _12904_/D _12900_/X VGND VGND VPWR VPWR _12901_/X sky130_fd_sc_hd__o22a_1
X_13881_ _13877_/X _13878_/X _13879_/X _13880_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13881_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15620_ _15621_/CLK _15620_/D VGND VGND VPWR VPWR pc[15] sky130_fd_sc_hd__dfxtp_2
XFILLER_36_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12832_ _12828_/X _12243_/X _12829_/X _12831_/X VGND VGND VPWR VPWR _12832_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_46_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15551_ _15591_/CLK _15551_/D VGND VGND VPWR VPWR _15551_/Q sky130_fd_sc_hd__dfxtp_1
X_12763_ _12763_/A VGND VGND VPWR VPWR _12763_/X sky130_fd_sc_hd__buf_1
X_14502_ _11676_/X _14502_/D VGND VGND VPWR VPWR _14502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11714_ _11723_/A VGND VGND VPWR VPWR _11714_/X sky130_fd_sc_hd__buf_1
X_15482_ _15509_/CLK _15482_/D VGND VGND VPWR VPWR wdata[8] sky130_fd_sc_hd__dfxtp_2
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12694_/A VGND VGND VPWR VPWR _12703_/B sky130_fd_sc_hd__buf_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _11917_/X _14433_/D VGND VGND VPWR VPWR _14433_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11647_/A VGND VGND VPWR VPWR _11645_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14364_ _15663_/CLK pc[25] VGND VGND VPWR VPWR _14364_/Q sky130_fd_sc_hd__dfxtp_1
X_11576_ _11576_/A _11798_/B VGND VGND VPWR VPWR _11589_/A sky130_fd_sc_hd__or2_2
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13315_ _12838_/X _12211_/X _13418_/S VGND VGND VPWR VPWR _13315_/X sky130_fd_sc_hd__mux2_1
X_10527_ _10536_/A VGND VGND VPWR VPWR _10527_/X sky130_fd_sc_hd__buf_1
X_14295_ _15510_/CLK _15462_/Q VGND VGND VPWR VPWR _14295_/Q sky130_fd_sc_hd__dfxtp_1
X_13246_ _13247_/X _13259_/X _13415_/S VGND VGND VPWR VPWR _13246_/X sky130_fd_sc_hd__mux2_1
X_10458_ _10460_/A VGND VGND VPWR VPWR _10458_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10389_ _10389_/A VGND VGND VPWR VPWR _10389_/X sky130_fd_sc_hd__buf_1
X_13177_ _12435_/X _12415_/X _13418_/S VGND VGND VPWR VPWR _13177_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12128_ _12128_/A VGND VGND VPWR VPWR _12148_/A sky130_fd_sc_hd__buf_1
XFILLER_123_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12059_ _12333_/B _12059_/B VGND VGND VPWR VPWR _12448_/A sky130_fd_sc_hd__or2_2
XFILLER_78_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09270_ _09278_/A VGND VGND VPWR VPWR _09270_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08221_ _08925_/A _09294_/B _11574_/C VGND VGND VPWR VPWR _08550_/B sky130_fd_sc_hd__or3_1
XFILLER_21_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08152_ _08182_/A VGND VGND VPWR VPWR _08173_/A sky130_fd_sc_hd__buf_2
XFILLER_147_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08083_ _14307_/Q VGND VGND VPWR VPWR _08084_/A sky130_fd_sc_hd__buf_1
XFILLER_107_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08985_ _08994_/A VGND VGND VPWR VPWR _08985_/X sky130_fd_sc_hd__buf_1
XFILLER_102_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07936_ _07936_/A VGND VGND VPWR VPWR _07936_/X sky130_fd_sc_hd__buf_1
XFILLER_87_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07867_ _07867_/A VGND VGND VPWR VPWR _07867_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09606_ _10745_/A VGND VGND VPWR VPWR _10363_/A sky130_fd_sc_hd__buf_1
XFILLER_84_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07798_ _07798_/A _07798_/B VGND VGND VPWR VPWR _07798_/X sky130_fd_sc_hd__or2_1
XFILLER_56_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09537_ _09551_/A VGND VGND VPWR VPWR _09537_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ _15059_/Q _09466_/X _09224_/X _09467_/X VGND VGND VPWR VPWR _15059_/D sky130_fd_sc_hd__a22o_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08419_ _10727_/A VGND VGND VPWR VPWR _09206_/A sky130_fd_sc_hd__buf_1
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09399_ _15078_/Q _09395_/X _09279_/X _09396_/X VGND VGND VPWR VPWR _15078_/D sky130_fd_sc_hd__a22o_1
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11430_ _11430_/A VGND VGND VPWR VPWR _11430_/X sky130_fd_sc_hd__buf_1
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11361_ _14583_/Q _11354_/X _11116_/X _11355_/X VGND VGND VPWR VPWR _14583_/D sky130_fd_sc_hd__a22o_1
X_13100_ _15646_/Q data_address[11] _15667_/Q VGND VGND VPWR VPWR _13100_/X sky130_fd_sc_hd__mux2_1
X_10312_ _10392_/A VGND VGND VPWR VPWR _10339_/A sky130_fd_sc_hd__buf_2
XFILLER_152_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11292_ _11301_/A VGND VGND VPWR VPWR _11299_/A sky130_fd_sc_hd__buf_1
X_14080_ _14968_/Q _15064_/Q _15032_/Q _15096_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14080_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10243_ _14866_/Q _10237_/X _10003_/X _10238_/X VGND VGND VPWR VPWR _14866_/D sky130_fd_sc_hd__a22o_1
X_13031_ wdata[4] rdata[4] _13058_/S VGND VGND VPWR VPWR _14308_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10174_ _10240_/A VGND VGND VPWR VPWR _10201_/A sky130_fd_sc_hd__buf_2
XFILLER_121_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14982_ _09800_/X _14982_/D VGND VGND VPWR VPWR _14982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13933_ _14662_/Q _15238_/Q _14726_/Q _14694_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13933_/X sky130_fd_sc_hd__mux4_2
XFILLER_75_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13864_ _15181_/Q _15149_/Q _14765_/Q _14797_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13864_/X sky130_fd_sc_hd__mux4_1
X_15603_ _15604_/CLK _15603_/D VGND VGND VPWR VPWR _15603_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ _12815_/A VGND VGND VPWR VPWR _12926_/A sky130_fd_sc_hd__buf_1
XFILLER_62_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13795_ _15124_/Q _15348_/Q _15316_/Q _15284_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13795_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15534_ _15566_/CLK _15534_/D VGND VGND VPWR VPWR _15534_/Q sky130_fd_sc_hd__dfxtp_1
X_12746_ _12746_/A VGND VGND VPWR VPWR _12746_/X sky130_fd_sc_hd__buf_1
XFILLER_43_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15465_ _15510_/CLK _15465_/D VGND VGND VPWR VPWR _15465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12677_ _12789_/A VGND VGND VPWR VPWR _12677_/X sky130_fd_sc_hd__buf_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ _11975_/X _14416_/D VGND VGND VPWR VPWR _14416_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11628_ _11628_/A VGND VGND VPWR VPWR _11628_/X sky130_fd_sc_hd__clkbuf_1
X_15396_ _08093_/X _15396_/D VGND VGND VPWR VPWR _15396_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14347_ _15621_/CLK pc[8] VGND VGND VPWR VPWR _14347_/Q sky130_fd_sc_hd__dfxtp_1
X_11559_ _11559_/A VGND VGND VPWR VPWR _11755_/A sky130_fd_sc_hd__buf_1
XFILLER_144_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14278_ _14500_/Q _14468_/Q _14436_/Q _14404_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14278_/X sky130_fd_sc_hd__mux4_2
Xrepeater5 _13649_/S VGND VGND VPWR VPWR _13641_/S sky130_fd_sc_hd__buf_6
X_13229_ _13228_/X _12884_/X _15565_/Q VGND VGND VPWR VPWR _13229_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08770_ _08770_/A VGND VGND VPWR VPWR _08770_/X sky130_fd_sc_hd__clkbuf_2
X_07721_ _07720_/A _07660_/A _07720_/Y VGND VGND VPWR VPWR _07722_/A sky130_fd_sc_hd__a21oi_2
XFILLER_84_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07652_ _07652_/A VGND VGND VPWR VPWR _07653_/A sky130_fd_sc_hd__buf_1
XFILLER_38_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07583_ _07585_/A _13079_/X VGND VGND VPWR VPWR _15494_/D sky130_fd_sc_hd__and2_1
XFILLER_81_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09322_ _09508_/A VGND VGND VPWR VPWR _09383_/A sky130_fd_sc_hd__buf_1
X_09253_ _15117_/Q _09249_/X _09250_/X _09252_/X VGND VGND VPWR VPWR _15117_/D sky130_fd_sc_hd__a22o_1
X_08204_ _08204_/A VGND VGND VPWR VPWR _08204_/X sky130_fd_sc_hd__buf_1
X_09184_ _09184_/A VGND VGND VPWR VPWR _09184_/X sky130_fd_sc_hd__buf_1
XFILLER_119_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08135_ _08144_/A VGND VGND VPWR VPWR _08135_/X sky130_fd_sc_hd__buf_1
XFILLER_146_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08066_ _15402_/Q _08062_/X _08064_/X _08065_/X VGND VGND VPWR VPWR _15402_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08968_ _08968_/A VGND VGND VPWR VPWR _08968_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07919_ _14297_/Q VGND VGND VPWR VPWR _07919_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08899_ _08921_/A VGND VGND VPWR VPWR _08908_/A sky130_fd_sc_hd__buf_1
X_10930_ _14696_/Q _10924_/X _10809_/X _10925_/X VGND VGND VPWR VPWR _14696_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10861_ _14717_/Q _10853_/X _10698_/X _10856_/X VGND VGND VPWR VPWR _14717_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12600_ _12739_/A VGND VGND VPWR VPWR _12600_/X sky130_fd_sc_hd__buf_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13580_ _14116_/X _14121_/X _13648_/S VGND VGND VPWR VPWR _13580_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10792_ _10802_/A VGND VGND VPWR VPWR _10792_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12531_ _12524_/A _12522_/A _15592_/Q _15560_/Q VGND VGND VPWR VPWR _12951_/C sky130_fd_sc_hd__o22a_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15250_ _08727_/X _15250_/D VGND VGND VPWR VPWR _15250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12462_ _12466_/A VGND VGND VPWR VPWR _12509_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14201_ _14197_/X _14198_/X _14199_/X _14200_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14201_/X sky130_fd_sc_hd__mux4_2
X_11413_ _11413_/A VGND VGND VPWR VPWR _11413_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15181_ _09004_/X _15181_/D VGND VGND VPWR VPWR _15181_/Q sky130_fd_sc_hd__dfxtp_1
X_12393_ _12388_/X _12392_/B _12401_/A VGND VGND VPWR VPWR _12394_/A sky130_fd_sc_hd__a21oi_4
XFILLER_126_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14132_ _15218_/Q _14546_/Q _14994_/Q _15410_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14132_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11344_ _11355_/A VGND VGND VPWR VPWR _11344_/X sky130_fd_sc_hd__buf_1
XFILLER_137_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14063_ _14681_/Q _15257_/Q _14745_/Q _14713_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14063_/X sky130_fd_sc_hd__mux4_2
X_11275_ _14608_/Q _11273_/X _11148_/X _11274_/X VGND VGND VPWR VPWR _14608_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13014_ _14358_/Q VGND VGND VPWR VPWR _13014_/Y sky130_fd_sc_hd__inv_2
X_10226_ _10256_/A VGND VGND VPWR VPWR _10247_/A sky130_fd_sc_hd__buf_2
XFILLER_67_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10157_ _10166_/A VGND VGND VPWR VPWR _10157_/X sky130_fd_sc_hd__buf_1
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14965_ _09863_/X _14965_/D VGND VGND VPWR VPWR _14965_/Q sky130_fd_sc_hd__dfxtp_1
X_10088_ _10148_/A VGND VGND VPWR VPWR _10107_/A sky130_fd_sc_hd__buf_2
XFILLER_63_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13916_ _13912_/X _13913_/X _13914_/X _13915_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13916_/X sky130_fd_sc_hd__mux4_2
XFILLER_75_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14896_ _10135_/X _14896_/D VGND VGND VPWR VPWR _14896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13847_ _14639_/Q _14607_/Q _14575_/Q _15375_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13847_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13778_ _14518_/Q _14486_/Q _14454_/Q _14422_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13778_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15517_ _15517_/CLK _15517_/D VGND VGND VPWR VPWR _15517_/Q sky130_fd_sc_hd__dfxtp_1
X_12729_ _12724_/X _12172_/X _12472_/X _12728_/X VGND VGND VPWR VPWR _12729_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_31_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15448_ _15669_/CLK _15448_/D VGND VGND VPWR VPWR data_address[21] sky130_fd_sc_hd__dfxtp_2
XFILLER_90_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15379_ _08163_/X _15379_/D VGND VGND VPWR VPWR _15379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09940_ _09949_/A VGND VGND VPWR VPWR _09940_/X sky130_fd_sc_hd__clkbuf_1
X_09871_ _09880_/A VGND VGND VPWR VPWR _09876_/A sky130_fd_sc_hd__buf_1
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08822_ _09192_/A VGND VGND VPWR VPWR _08822_/X sky130_fd_sc_hd__buf_1
XFILLER_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08753_ _08762_/A VGND VGND VPWR VPWR _08753_/X sky130_fd_sc_hd__buf_1
X_07704_ _07701_/X _13133_/X _07701_/X _13133_/X VGND VGND VPWR VPWR _07705_/A sky130_fd_sc_hd__a2bb2o_1
X_08684_ _09000_/A VGND VGND VPWR VPWR _08897_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07635_ _07635_/A _12030_/C VGND VGND VPWR VPWR _15464_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07566_ _07557_/X _07560_/Y _07562_/X _07565_/X VGND VGND VPWR VPWR _15506_/D sky130_fd_sc_hd__o211a_1
XFILLER_34_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09305_ _09305_/A VGND VGND VPWR VPWR _09305_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07497_ _07500_/A _07497_/B VGND VGND VPWR VPWR _15523_/D sky130_fd_sc_hd__nor2_1
X_09236_ _09236_/A VGND VGND VPWR VPWR _09236_/X sky130_fd_sc_hd__buf_1
XFILLER_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09167_ _09167_/A VGND VGND VPWR VPWR _09248_/A sky130_fd_sc_hd__buf_2
XFILLER_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08118_ _08118_/A VGND VGND VPWR VPWR _08129_/A sky130_fd_sc_hd__buf_1
XFILLER_119_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09098_ _09202_/A VGND VGND VPWR VPWR _09161_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08049_ _08049_/A VGND VGND VPWR VPWR _08080_/A sky130_fd_sc_hd__buf_1
XFILLER_122_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11060_ _11070_/A VGND VGND VPWR VPWR _11060_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10011_ _10011_/A VGND VGND VPWR VPWR _10011_/X sky130_fd_sc_hd__buf_1
XFILLER_89_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14750_ _10689_/X _14750_/D VGND VGND VPWR VPWR _14750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11962_ _11962_/A VGND VGND VPWR VPWR _11962_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13701_ _13697_/X _13698_/X _13699_/X _13700_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13701_/X sky130_fd_sc_hd__mux4_1
X_10913_ _10913_/A VGND VGND VPWR VPWR _10936_/A sky130_fd_sc_hd__buf_1
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14681_ _10984_/X _14681_/D VGND VGND VPWR VPWR _14681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11893_ _14440_/Q _11886_/X _08074_/A _11887_/X VGND VGND VPWR VPWR _14440_/D sky130_fd_sc_hd__a22o_1
X_13632_ _14246_/X _14251_/X _13648_/S VGND VGND VPWR VPWR _13632_/X sky130_fd_sc_hd__mux2_2
X_10844_ _14722_/Q _10840_/X _10665_/X _10843_/X VGND VGND VPWR VPWR _14722_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13563_ _13562_/X _13081_/X _14337_/Q VGND VGND VPWR VPWR _13563_/X sky130_fd_sc_hd__mux2_1
X_10775_ _10775_/A VGND VGND VPWR VPWR _11523_/A sky130_fd_sc_hd__clkbuf_2
X_15302_ _08526_/X _15302_/D VGND VGND VPWR VPWR _15302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12514_ _12513_/A _12513_/B _12512_/X _12513_/Y VGND VGND VPWR VPWR _12514_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13494_ _13876_/X _13881_/X _13521_/S VGND VGND VPWR VPWR _13494_/X sky130_fd_sc_hd__mux2_2
X_15233_ _08788_/X _15233_/D VGND VGND VPWR VPWR _15233_/Q sky130_fd_sc_hd__dfxtp_1
X_12445_ _12670_/A VGND VGND VPWR VPWR _12593_/A sky130_fd_sc_hd__clkbuf_2
X_15164_ _09064_/X _15164_/D VGND VGND VPWR VPWR _15164_/Q sky130_fd_sc_hd__dfxtp_1
X_12376_ _12400_/B _13345_/X VGND VGND VPWR VPWR _12376_/X sky130_fd_sc_hd__or2_2
X_14115_ _15124_/Q _15348_/Q _15316_/Q _15284_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14115_/X sky130_fd_sc_hd__mux4_1
X_11327_ _11329_/A VGND VGND VPWR VPWR _11327_/X sky130_fd_sc_hd__clkbuf_1
X_15095_ _09340_/X _15095_/D VGND VGND VPWR VPWR _15095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14046_ _14042_/X _14043_/X _14044_/X _14045_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14046_/X sky130_fd_sc_hd__mux4_2
X_11258_ _11260_/A VGND VGND VPWR VPWR _11258_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10209_ _14876_/Q _10207_/X _09958_/X _10208_/X VGND VGND VPWR VPWR _14876_/D sky130_fd_sc_hd__a22o_1
X_11189_ _14631_/Q _11186_/X _11187_/X _11188_/X VGND VGND VPWR VPWR _14631_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14948_ _09915_/X _14948_/D VGND VGND VPWR VPWR _14948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14879_ _10193_/X _14879_/D VGND VGND VPWR VPWR _14879_/Q sky130_fd_sc_hd__dfxtp_1
X_07420_ _07420_/A VGND VGND VPWR VPWR _07429_/A sky130_fd_sc_hd__buf_1
XFILLER_63_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07351_ _07497_/B _07339_/X _07498_/B _07341_/X VGND VGND VPWR VPWR _07353_/B sky130_fd_sc_hd__o22a_2
XFILLER_50_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07282_ _07282_/A _07282_/B VGND VGND VPWR VPWR _15613_/D sky130_fd_sc_hd__nor2_1
XFILLER_148_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09021_ _09021_/A VGND VGND VPWR VPWR _09021_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09923_ _09923_/A _09923_/B _14301_/Q VGND VGND VPWR VPWR _10294_/B sky130_fd_sc_hd__or3_1
XFILLER_120_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09854_ _09854_/A VGND VGND VPWR VPWR _09854_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08805_ _09176_/A VGND VGND VPWR VPWR _08805_/X sky130_fd_sc_hd__buf_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09785_ _09785_/A VGND VGND VPWR VPWR _09792_/A sky130_fd_sc_hd__buf_1
XFILLER_85_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08736_ _08740_/A VGND VGND VPWR VPWR _08736_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_107 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_118 rdata[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08667_ _08677_/A VGND VGND VPWR VPWR _08680_/A sky130_fd_sc_hd__inv_2
XANTENNA_129 rdata[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07618_ _12036_/A VGND VGND VPWR VPWR _07619_/B sky130_fd_sc_hd__buf_1
XFILLER_14_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08598_ _08628_/A VGND VGND VPWR VPWR _08618_/A sky130_fd_sc_hd__clkbuf_2
X_07549_ _15515_/Q VGND VGND VPWR VPWR _07632_/B sky130_fd_sc_hd__inv_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10560_ _14784_/Q _10550_/X _10308_/X _10553_/X VGND VGND VPWR VPWR _14784_/D sky130_fd_sc_hd__a22o_1
X_09219_ _09227_/A VGND VGND VPWR VPWR _09219_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10491_ _14804_/Q _10484_/X _10363_/X _10486_/X VGND VGND VPWR VPWR _14804_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12230_ _12230_/A _12230_/B VGND VGND VPWR VPWR _12230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12161_ _12709_/A _12160_/B _12690_/A VGND VGND VPWR VPWR _12689_/A sky130_fd_sc_hd__a21boi_4
XFILLER_146_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11112_ _11479_/A VGND VGND VPWR VPWR _11112_/X sky130_fd_sc_hd__buf_1
XFILLER_146_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12092_ _12092_/A VGND VGND VPWR VPWR _12092_/X sky130_fd_sc_hd__buf_1
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11043_ _11045_/A VGND VGND VPWR VPWR _11043_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14802_ _10499_/X _14802_/D VGND VGND VPWR VPWR _14802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12994_ _15506_/D VGND VGND VPWR VPWR _15672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14733_ _10778_/X _14733_/D VGND VGND VPWR VPWR _14733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11945_ _11951_/A VGND VGND VPWR VPWR _11945_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14664_ _11043_/X _14664_/D VGND VGND VPWR VPWR _14664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11876_ _11876_/A VGND VGND VPWR VPWR _11896_/A sky130_fd_sc_hd__clkbuf_2
X_13615_ _13614_/X _13068_/X _14337_/Q VGND VGND VPWR VPWR _13615_/X sky130_fd_sc_hd__mux2_1
X_10827_ _10827_/A VGND VGND VPWR VPWR _11567_/A sky130_fd_sc_hd__buf_1
X_14595_ _11314_/X _14595_/D VGND VGND VPWR VPWR _14595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13546_ _13545_/X _14330_/D _15506_/Q VGND VGND VPWR VPWR _13546_/X sky130_fd_sc_hd__mux2_1
X_10758_ _10773_/A VGND VGND VPWR VPWR _10769_/A sky130_fd_sc_hd__buf_1
XFILLER_9_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13477_ _13476_/X rdata[15] _13516_/S VGND VGND VPWR VPWR _13477_/X sky130_fd_sc_hd__mux2_1
X_10689_ _10689_/A VGND VGND VPWR VPWR _10689_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15216_ _08863_/X _15216_/D VGND VGND VPWR VPWR _15216_/Q sky130_fd_sc_hd__dfxtp_1
X_12428_ _12428_/A VGND VGND VPWR VPWR _12428_/X sky130_fd_sc_hd__buf_2
X_15147_ _09123_/X _15147_/D VGND VGND VPWR VPWR _15147_/Q sky130_fd_sc_hd__dfxtp_1
X_12359_ _15554_/Q VGND VGND VPWR VPWR _12359_/X sky130_fd_sc_hd__buf_1
XFILLER_99_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15078_ _09398_/X _15078_/D VGND VGND VPWR VPWR _15078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14029_ _14845_/Q _14877_/Q _14909_/Q _14941_/Q _14060_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14029_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09570_ _15035_/Q _09562_/X _09569_/X _09565_/X VGND VGND VPWR VPWR _15035_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08521_ _14308_/Q VGND VGND VPWR VPWR _10813_/A sky130_fd_sc_hd__buf_1
XFILLER_35_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08452_ _14319_/Q VGND VGND VPWR VPWR _10755_/A sky130_fd_sc_hd__buf_1
XFILLER_50_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07403_ _07403_/A VGND VGND VPWR VPWR _07406_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_51_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08383_ _10697_/A VGND VGND VPWR VPWR _09180_/A sky130_fd_sc_hd__clkbuf_2
X_07334_ _14391_/Q VGND VGND VPWR VPWR _07494_/B sky130_fd_sc_hd__inv_2
XFILLER_50_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07265_ _07265_/A _07265_/B VGND VGND VPWR VPWR _15625_/D sky130_fd_sc_hd__nor2_4
X_09004_ _09012_/A VGND VGND VPWR VPWR _09004_/X sky130_fd_sc_hd__clkbuf_1
X_07196_ _07256_/B _07175_/B _07188_/X _07194_/Y VGND VGND VPWR VPWR _15661_/D sky130_fd_sc_hd__a211oi_4
XFILLER_129_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09906_ _09906_/A VGND VGND VPWR VPWR _09906_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09837_ _09846_/A VGND VGND VPWR VPWR _09837_/X sky130_fd_sc_hd__buf_1
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09768_ _09768_/A VGND VGND VPWR VPWR _09768_/X sky130_fd_sc_hd__buf_1
XFILLER_132_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08719_ _15253_/Q _08712_/X _08434_/X _08714_/X VGND VGND VPWR VPWR _15253_/D sky130_fd_sc_hd__a22o_1
X_09699_ _09709_/A VGND VGND VPWR VPWR _09699_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11730_ _14487_/Q _11722_/X _11484_/X _11723_/X VGND VGND VPWR VPWR _14487_/D sky130_fd_sc_hd__a22o_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11661_ _11725_/A VGND VGND VPWR VPWR _11680_/A sky130_fd_sc_hd__clkbuf_2
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _12329_/X _12395_/A _13418_/S VGND VGND VPWR VPWR _13400_/X sky130_fd_sc_hd__mux2_1
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10612_ _14770_/Q _10607_/X _10371_/X _10608_/X VGND VGND VPWR VPWR _14770_/D sky130_fd_sc_hd__a22o_1
X_14380_ _15646_/CLK instruction[9] VGND VGND VPWR VPWR _14380_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11592_ _11592_/A VGND VGND VPWR VPWR _11653_/A sky130_fd_sc_hd__buf_2
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ _13333_/X _13332_/X _13408_/S VGND VGND VPWR VPWR _13331_/X sky130_fd_sc_hd__mux2_1
X_10543_ _10547_/A VGND VGND VPWR VPWR _10543_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13262_ _13263_/X _12860_/B _13393_/S VGND VGND VPWR VPWR _13262_/X sky130_fd_sc_hd__mux2_2
X_10474_ _10474_/A VGND VGND VPWR VPWR _10474_/X sky130_fd_sc_hd__buf_1
XFILLER_108_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15001_ _09735_/X _15001_/D VGND VGND VPWR VPWR _15001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12213_ _15564_/Q VGND VGND VPWR VPWR _12213_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13193_ _13196_/X _13216_/X _13408_/S VGND VGND VPWR VPWR _13193_/X sky130_fd_sc_hd__mux2_1
X_12144_ _12144_/A _12144_/B _12636_/A VGND VGND VPWR VPWR _12144_/X sky130_fd_sc_hd__or3b_4
X_12075_ _12577_/A _12075_/B VGND VGND VPWR VPWR _12076_/A sky130_fd_sc_hd__or2_1
X_11026_ _11026_/A VGND VGND VPWR VPWR _11047_/A sky130_fd_sc_hd__buf_1
XFILLER_110_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12977_ _12977_/A VGND VGND VPWR VPWR _12984_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14716_ _10863_/X _14716_/D VGND VGND VPWR VPWR _14716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11928_ _11947_/A VGND VGND VPWR VPWR _11928_/X sky130_fd_sc_hd__buf_1
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14647_ _11115_/X _14647_/D VGND VGND VPWR VPWR _14647_/Q sky130_fd_sc_hd__dfxtp_1
X_11859_ _11859_/A VGND VGND VPWR VPWR _11859_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_18 data_address[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ _11379_/X _14578_/D VGND VGND VPWR VPWR _14578_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_29 data_address[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13529_ _13528_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13529_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07952_ _07952_/A VGND VGND VPWR VPWR _08049_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07883_ _07878_/A _07878_/B _07882_/X _07878_/Y VGND VGND VPWR VPWR _15437_/D sky130_fd_sc_hd__o211a_1
XFILLER_96_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09622_ _10375_/A VGND VGND VPWR VPWR _09622_/X sky130_fd_sc_hd__buf_1
XFILLER_110_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09553_ _10320_/A VGND VGND VPWR VPWR _09553_/X sky130_fd_sc_hd__buf_1
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08504_ _10798_/A VGND VGND VPWR VPWR _09263_/A sky130_fd_sc_hd__buf_1
X_09484_ _09484_/A VGND VGND VPWR VPWR _09484_/X sky130_fd_sc_hd__clkbuf_1
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08435_ _15317_/Q _08424_/X _08434_/X _08429_/X VGND VGND VPWR VPWR _15317_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ _08405_/A VGND VGND VPWR VPWR _08366_/X sky130_fd_sc_hd__buf_1
XFILLER_20_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07317_ _07321_/B _07321_/C _07513_/B VGND VGND VPWR VPWR _07338_/A sky130_fd_sc_hd__or3_1
X_08297_ _08583_/A VGND VGND VPWR VPWR _08379_/A sky130_fd_sc_hd__buf_2
XFILLER_20_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07248_ _07274_/A VGND VGND VPWR VPWR _07257_/A sky130_fd_sc_hd__buf_1
XFILLER_127_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07179_ _07251_/B _07179_/B VGND VGND VPWR VPWR _07180_/A sky130_fd_sc_hd__or2_1
XFILLER_105_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10190_ _14881_/Q _10183_/X _09934_/X _10186_/X VGND VGND VPWR VPWR _14881_/D sky130_fd_sc_hd__a22o_1
XFILLER_132_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12900_ _12386_/Y _12379_/B _12904_/B _12899_/X VGND VGND VPWR VPWR _12900_/X sky130_fd_sc_hd__o22a_1
XFILLER_101_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13880_ _14956_/Q _15052_/Q _15020_/Q _15084_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13880_/X sky130_fd_sc_hd__mux4_2
XFILLER_46_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12831_ _12820_/X _12825_/X _12830_/X VGND VGND VPWR VPWR _12831_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15550_ _15591_/CLK _15550_/D VGND VGND VPWR VPWR _15550_/Q sky130_fd_sc_hd__dfxtp_1
X_12762_ _12762_/A VGND VGND VPWR VPWR _12762_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_15_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14501_ _11678_/X _14501_/D VGND VGND VPWR VPWR _14501_/Q sky130_fd_sc_hd__dfxtp_1
X_11713_ _11722_/A VGND VGND VPWR VPWR _11713_/X sky130_fd_sc_hd__buf_1
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15481_ _15509_/CLK _15481_/D VGND VGND VPWR VPWR wdata[7] sky130_fd_sc_hd__dfxtp_2
XFILLER_70_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12693_ _12693_/A VGND VGND VPWR VPWR _12703_/A sky130_fd_sc_hd__buf_2
XFILLER_70_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _11919_/X _14432_/D VGND VGND VPWR VPWR _14432_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _14512_/Q _11642_/X _11514_/X _11643_/X VGND VGND VPWR VPWR _14512_/D sky130_fd_sc_hd__a22o_1
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ _15663_/CLK pc[24] VGND VGND VPWR VPWR _14363_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11575_ _11910_/B VGND VGND VPWR VPWR _11798_/B sky130_fd_sc_hd__clkbuf_1
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13314_ _13315_/X _13339_/X _13415_/S VGND VGND VPWR VPWR _13314_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10526_ _10535_/A VGND VGND VPWR VPWR _10526_/X sky130_fd_sc_hd__buf_1
X_14294_ _15510_/CLK _15461_/Q VGND VGND VPWR VPWR _14294_/Q sky130_fd_sc_hd__dfxtp_1
X_13245_ _13246_/X _13270_/X _13408_/S VGND VGND VPWR VPWR _13245_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10457_ _14815_/Q _10453_/X _10314_/X _10456_/X VGND VGND VPWR VPWR _14815_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13176_ _13175_/X _13256_/X _15565_/Q VGND VGND VPWR VPWR _13176_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10388_ _10398_/A VGND VGND VPWR VPWR _10388_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12127_ _15577_/Q VGND VGND VPWR VPWR _12675_/A sky130_fd_sc_hd__inv_2
XFILLER_151_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12058_ _12316_/B _12307_/B VGND VGND VPWR VPWR _12059_/B sky130_fd_sc_hd__or2_1
X_11009_ _11018_/A VGND VGND VPWR VPWR _11014_/A sky130_fd_sc_hd__buf_1
XFILLER_92_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_opt_2_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR clkbuf_opt_2_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08220_ _08662_/C VGND VGND VPWR VPWR _11574_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_60_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08151_ _08159_/A VGND VGND VPWR VPWR _08151_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08082_ _08082_/A VGND VGND VPWR VPWR _08082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08984_ _08993_/A VGND VGND VPWR VPWR _08984_/X sky130_fd_sc_hd__buf_1
X_07935_ _14334_/Q VGND VGND VPWR VPWR _07936_/A sky130_fd_sc_hd__buf_1
XFILLER_29_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07866_ _07848_/X _07709_/X _07872_/B VGND VGND VPWR VPWR _07867_/A sky130_fd_sc_hd__o21ai_2
XFILLER_110_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09605_ _09615_/A VGND VGND VPWR VPWR _09605_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07797_ _07789_/A _07789_/B _07796_/X _07789_/Y VGND VGND VPWR VPWR _15457_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09536_ _09536_/A VGND VGND VPWR VPWR _09551_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09467_ _09476_/A VGND VGND VPWR VPWR _09467_/X sky130_fd_sc_hd__buf_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08418_ _14324_/Q VGND VGND VPWR VPWR _10727_/A sky130_fd_sc_hd__buf_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09398_ _09400_/A VGND VGND VPWR VPWR _09398_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08349_ _08370_/A VGND VGND VPWR VPWR _08350_/A sky130_fd_sc_hd__buf_1
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11360_ _11362_/A VGND VGND VPWR VPWR _11360_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10311_ _10311_/A VGND VGND VPWR VPWR _10392_/A sky130_fd_sc_hd__buf_2
XFILLER_138_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11291_ _14603_/Q _11284_/X _11170_/X _11286_/X VGND VGND VPWR VPWR _14603_/D sky130_fd_sc_hd__a22o_1
X_13030_ wdata[3] rdata[3] _13058_/S VGND VGND VPWR VPWR _14307_/D sky130_fd_sc_hd__mux2_1
X_10242_ _10246_/A VGND VGND VPWR VPWR _10242_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10173_ _10173_/A VGND VGND VPWR VPWR _10240_/A sky130_fd_sc_hd__buf_1
XFILLER_133_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14981_ _09802_/X _14981_/D VGND VGND VPWR VPWR _14981_/Q sky130_fd_sc_hd__dfxtp_1
X_13932_ _15206_/Q _14534_/Q _14982_/Q _15398_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13932_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13863_ _14669_/Q _15245_/Q _14733_/Q _14701_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13863_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15602_ _15667_/CLK _15602_/D VGND VGND VPWR VPWR _15602_/Q sky130_fd_sc_hd__dfxtp_1
X_12814_ _12745_/X _12804_/Y _12809_/Y _12813_/X VGND VGND VPWR VPWR _12814_/Y sky130_fd_sc_hd__o211ai_1
X_13794_ _15188_/Q _15156_/Q _14772_/Q _14804_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13794_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12745_ _12745_/A VGND VGND VPWR VPWR _12745_/X sky130_fd_sc_hd__buf_1
X_15533_ _15578_/CLK _15533_/D VGND VGND VPWR VPWR _15533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15464_ _15604_/CLK _15464_/D VGND VGND VPWR VPWR _15464_/Q sky130_fd_sc_hd__dfxtp_1
X_12676_ _12676_/A VGND VGND VPWR VPWR _12676_/X sky130_fd_sc_hd__buf_1
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _11979_/X _14415_/D VGND VGND VPWR VPWR _14415_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _14517_/Q _11622_/X _11494_/X _11624_/X VGND VGND VPWR VPWR _14517_/D sky130_fd_sc_hd__a22o_1
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15395_ _08097_/X _15395_/D VGND VGND VPWR VPWR _15395_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ _15601_/CLK pc[7] VGND VGND VPWR VPWR _14346_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ _14534_/Q _11552_/X _11557_/X _11554_/X VGND VGND VPWR VPWR _14534_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10509_ _14799_/Q _10505_/X _10383_/X _10506_/X VGND VGND VPWR VPWR _14799_/D sky130_fd_sc_hd__a22o_1
XFILLER_128_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14277_ _14628_/Q _14596_/Q _14564_/Q _15364_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14277_/X sky130_fd_sc_hd__mux4_2
X_11489_ _11489_/A VGND VGND VPWR VPWR _11489_/X sky130_fd_sc_hd__buf_1
Xrepeater6 _13058_/S VGND VGND VPWR VPWR _13057_/S sky130_fd_sc_hd__buf_8
X_13228_ _13230_/X _13275_/X _15564_/Q VGND VGND VPWR VPWR _13228_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13159_ _13158_/X _13172_/X _15562_/Q VGND VGND VPWR VPWR _13159_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07720_ _07720_/A _15604_/Q VGND VGND VPWR VPWR _07720_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07651_ _07689_/A VGND VGND VPWR VPWR _07652_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_66_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07582_ _07582_/A VGND VGND VPWR VPWR _07585_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09321_ _09964_/A VGND VGND VPWR VPWR _09508_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_34_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09252_ _09276_/A VGND VGND VPWR VPWR _09252_/X sky130_fd_sc_hd__buf_1
XFILLER_33_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08203_ _08209_/A VGND VGND VPWR VPWR _08203_/X sky130_fd_sc_hd__clkbuf_1
X_09183_ _09195_/A VGND VGND VPWR VPWR _09183_/X sky130_fd_sc_hd__buf_1
X_08134_ _08143_/A VGND VGND VPWR VPWR _08134_/X sky130_fd_sc_hd__buf_1
XFILLER_146_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08065_ _08080_/A VGND VGND VPWR VPWR _08065_/X sky130_fd_sc_hd__buf_1
XFILLER_135_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08967_ _15192_/Q _08963_/X _08830_/X _08964_/X VGND VGND VPWR VPWR _15192_/D sky130_fd_sc_hd__a22o_1
X_07918_ _14300_/Q VGND VGND VPWR VPWR _08340_/B sky130_fd_sc_hd__inv_2
XFILLER_84_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08898_ _08970_/A VGND VGND VPWR VPWR _08921_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07849_ _07849_/A _07854_/A VGND VGND VPWR VPWR _07849_/X sky130_fd_sc_hd__or2_1
XFILLER_44_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10860_ _10860_/A VGND VGND VPWR VPWR _10860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09519_ _15043_/Q _09410_/A _09290_/X _09413_/A VGND VGND VPWR VPWR _15043_/D sky130_fd_sc_hd__a22o_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10791_ _10821_/A VGND VGND VPWR VPWR _10802_/A sky130_fd_sc_hd__buf_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _12530_/A VGND VGND VPWR VPWR _12530_/Y sky130_fd_sc_hd__inv_2
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12461_ _15558_/Q VGND VGND VPWR VPWR _12466_/A sky130_fd_sc_hd__inv_2
X_14200_ _14956_/Q _15052_/Q _15020_/Q _15084_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14200_/X sky130_fd_sc_hd__mux4_2
XFILLER_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11412_ _14568_/Q _11404_/X _11183_/X _11405_/X VGND VGND VPWR VPWR _14568_/D sky130_fd_sc_hd__a22o_1
X_15180_ _09010_/X _15180_/D VGND VGND VPWR VPWR _15180_/Q sky130_fd_sc_hd__dfxtp_1
X_12392_ _12392_/A _12392_/B VGND VGND VPWR VPWR _12401_/A sky130_fd_sc_hd__nor2_2
XFILLER_153_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14131_ _14127_/X _14128_/X _14129_/X _14130_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14131_/X sky130_fd_sc_hd__mux4_2
X_11343_ _11354_/A VGND VGND VPWR VPWR _11343_/X sky130_fd_sc_hd__buf_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14062_ _15225_/Q _14553_/Q _15001_/Q _15417_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14062_/X sky130_fd_sc_hd__mux4_1
X_11274_ _11274_/A VGND VGND VPWR VPWR _11274_/X sky130_fd_sc_hd__buf_1
XFILLER_4_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13013_ _14357_/Q VGND VGND VPWR VPWR _13013_/Y sky130_fd_sc_hd__inv_2
X_10225_ _10225_/A VGND VGND VPWR VPWR _10225_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10156_ _10162_/A VGND VGND VPWR VPWR _10156_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14964_ _09865_/X _14964_/D VGND VGND VPWR VPWR _14964_/Q sky130_fd_sc_hd__dfxtp_1
X_10087_ _10087_/A VGND VGND VPWR VPWR _10148_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13915_ _15112_/Q _15336_/Q _15304_/Q _15272_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13915_/X sky130_fd_sc_hd__mux4_1
X_14895_ _10139_/X _14895_/D VGND VGND VPWR VPWR _14895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13846_ _13842_/X _13843_/X _13844_/X _13845_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13846_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13777_ _14646_/Q _14614_/Q _14582_/Q _15382_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13777_/X sky130_fd_sc_hd__mux4_2
X_10989_ _10993_/A VGND VGND VPWR VPWR _10989_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_90_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15516_ _15521_/CLK _15516_/D VGND VGND VPWR VPWR _15516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12728_ _12730_/A _12730_/B _12727_/X VGND VGND VPWR VPWR _12728_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15447_ _15456_/CLK _15447_/D VGND VGND VPWR VPWR data_address[20] sky130_fd_sc_hd__dfxtp_2
X_12659_ _12535_/X _12641_/B _12651_/Y _12653_/X _12658_/X VGND VGND VPWR VPWR _12660_/A
+ sky130_fd_sc_hd__o311a_1
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15378_ _08167_/X _15378_/D VGND VGND VPWR VPWR _15378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14329_ _15502_/CLK _14329_/D VGND VGND VPWR VPWR _14329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09870_ _14963_/Q _09868_/X _09612_/X _09869_/X VGND VGND VPWR VPWR _14963_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08821_ _08829_/A VGND VGND VPWR VPWR _08821_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08752_ _08752_/A VGND VGND VPWR VPWR _08752_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07703_ _07854_/A _07852_/A VGND VGND VPWR VPWR _07703_/X sky130_fd_sc_hd__or2_1
XFILLER_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08683_ _15263_/Q _08679_/X _08369_/X _08682_/X VGND VGND VPWR VPWR _15263_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07634_ _07634_/A _07634_/B VGND VGND VPWR VPWR _15465_/D sky130_fd_sc_hd__nor2_1
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07565_ _07379_/A _07535_/Y _12571_/A _15468_/Q _07564_/X VGND VGND VPWR VPWR _07565_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09304_ _15105_/Q _09298_/X _09159_/X _09301_/X VGND VGND VPWR VPWR _15105_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07496_ _07496_/A VGND VGND VPWR VPWR _07500_/A sky130_fd_sc_hd__buf_1
X_09235_ _09235_/A VGND VGND VPWR VPWR _09235_/X sky130_fd_sc_hd__buf_1
XFILLER_139_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09166_ _09175_/A VGND VGND VPWR VPWR _09166_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08117_ _15392_/Q _08109_/X _07944_/X _08112_/X VGND VGND VPWR VPWR _15392_/D sky130_fd_sc_hd__a22o_1
X_09097_ _15155_/Q _09095_/X _08852_/X _09096_/X VGND VGND VPWR VPWR _15155_/D sky130_fd_sc_hd__a22o_1
XFILLER_107_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08048_ _08048_/A VGND VGND VPWR VPWR _08048_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10010_ _10015_/A VGND VGND VPWR VPWR _10010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09999_ _10367_/A VGND VGND VPWR VPWR _09999_/X sky130_fd_sc_hd__buf_1
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11961_ _14421_/Q _11956_/X _08006_/A _11958_/X VGND VGND VPWR VPWR _14421_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10912_ _10920_/A VGND VGND VPWR VPWR _10912_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13700_ _14974_/Q _15070_/Q _15038_/Q _15102_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13700_/X sky130_fd_sc_hd__mux4_2
X_14680_ _10989_/X _14680_/D VGND VGND VPWR VPWR _14680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11892_ _11898_/A VGND VGND VPWR VPWR _11892_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13631_ _13630_/X _13064_/X _14337_/Q VGND VGND VPWR VPWR _13631_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10843_ _10843_/A VGND VGND VPWR VPWR _10843_/X sky130_fd_sc_hd__buf_1
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13562_ _13561_/X _14326_/D _15506_/Q VGND VGND VPWR VPWR _13562_/X sky130_fd_sc_hd__mux2_2
X_10774_ _10786_/A VGND VGND VPWR VPWR _10774_/X sky130_fd_sc_hd__clkbuf_1
X_12513_ _12513_/A _12513_/B VGND VGND VPWR VPWR _12513_/Y sky130_fd_sc_hd__nand2_1
X_15301_ _08532_/X _15301_/D VGND VGND VPWR VPWR _15301_/Q sky130_fd_sc_hd__dfxtp_1
X_13493_ _13492_/X _13069_/X _14336_/Q VGND VGND VPWR VPWR _13493_/X sky130_fd_sc_hd__mux2_1
X_12444_ _15589_/Q _15557_/Q VGND VGND VPWR VPWR _12444_/Y sky130_fd_sc_hd__nor2_1
X_15232_ _08792_/X _15232_/D VGND VGND VPWR VPWR _15232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15163_ _09070_/X _15163_/D VGND VGND VPWR VPWR _15163_/Q sky130_fd_sc_hd__dfxtp_1
X_12375_ _12349_/X _12358_/X _12361_/Y _12366_/X _12374_/X VGND VGND VPWR VPWR _12375_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14114_ _15188_/Q _15156_/Q _14772_/Q _14804_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14114_/X sky130_fd_sc_hd__mux4_1
X_11326_ _14593_/Q _11319_/X _11071_/X _11322_/X VGND VGND VPWR VPWR _14593_/D sky130_fd_sc_hd__a22o_1
XFILLER_126_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15094_ _09343_/X _15094_/D VGND VGND VPWR VPWR _15094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14045_ _15131_/Q _15355_/Q _15323_/Q _15291_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14045_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11257_ _14614_/Q _11254_/X _11121_/X _11256_/X VGND VGND VPWR VPWR _14614_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10208_ _10218_/A VGND VGND VPWR VPWR _10208_/X sky130_fd_sc_hd__buf_1
X_11188_ _11188_/A VGND VGND VPWR VPWR _11188_/X sky130_fd_sc_hd__buf_1
XFILLER_121_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10139_ _10141_/A VGND VGND VPWR VPWR _10139_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14947_ _09919_/X _14947_/D VGND VGND VPWR VPWR _14947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14878_ _10202_/X _14878_/D VGND VGND VPWR VPWR _14878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13829_ _14833_/Q _14865_/Q _14897_/Q _14929_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13829_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07350_ _14388_/Q VGND VGND VPWR VPWR _07498_/B sky130_fd_sc_hd__inv_2
XFILLER_31_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07281_ _07282_/A _07281_/B VGND VGND VPWR VPWR _15614_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09020_ _15177_/Q _09016_/X _08895_/X _09017_/X VGND VGND VPWR VPWR _15177_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09922_ _09922_/A VGND VGND VPWR VPWR _10838_/A sky130_fd_sc_hd__buf_1
X_09853_ _14967_/Q _09846_/X _09589_/X _09847_/X VGND VGND VPWR VPWR _14967_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08804_ _08804_/A VGND VGND VPWR VPWR _08804_/X sky130_fd_sc_hd__clkbuf_1
X_09784_ _14987_/Q _09777_/X _09657_/X _09779_/X VGND VGND VPWR VPWR _14987_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08735_ _08735_/A VGND VGND VPWR VPWR _08740_/A sky130_fd_sc_hd__buf_1
XFILLER_73_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_108 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_119 rdata[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08666_ _08666_/A VGND VGND VPWR VPWR _08666_/X sky130_fd_sc_hd__buf_1
X_07617_ _07617_/A VGND VGND VPWR VPWR _12036_/A sky130_fd_sc_hd__buf_1
XFILLER_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08597_ _08617_/A VGND VGND VPWR VPWR _08597_/X sky130_fd_sc_hd__buf_1
XFILLER_81_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07548_ _07628_/B _13521_/S _07633_/B _07542_/A VGND VGND VPWR VPWR _07556_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07479_ _07483_/A VGND VGND VPWR VPWR _07482_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09218_ _09230_/A VGND VGND VPWR VPWR _09227_/A sky130_fd_sc_hd__buf_1
X_10490_ _10490_/A VGND VGND VPWR VPWR _10490_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09149_ _09158_/A VGND VGND VPWR VPWR _09149_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12160_ _12160_/A _12160_/B VGND VGND VPWR VPWR _12690_/A sky130_fd_sc_hd__or2_1
XFILLER_135_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11111_ _11111_/A VGND VGND VPWR VPWR _11111_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12091_ _15581_/Q VGND VGND VPWR VPWR _12091_/X sky130_fd_sc_hd__buf_1
X_11042_ _14665_/Q _11037_/X _10804_/X _11038_/X VGND VGND VPWR VPWR _14665_/D sky130_fd_sc_hd__a22o_1
XFILLER_131_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14801_ _10501_/X _14801_/D VGND VGND VPWR VPWR _14801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12993_ _12993_/A _12993_/B VGND VGND VPWR VPWR _12993_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14732_ _10786_/X _14732_/D VGND VGND VPWR VPWR _14732_/Q sky130_fd_sc_hd__dfxtp_1
X_11944_ _11964_/A VGND VGND VPWR VPWR _11951_/A sky130_fd_sc_hd__buf_1
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14663_ _11045_/X _14663_/D VGND VGND VPWR VPWR _14663_/Q sky130_fd_sc_hd__dfxtp_1
X_11875_ _11895_/A VGND VGND VPWR VPWR _11875_/X sky130_fd_sc_hd__buf_1
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13614_ _13613_/X _14313_/D _15506_/Q VGND VGND VPWR VPWR _13614_/X sky130_fd_sc_hd__mux2_1
X_10826_ _10830_/A VGND VGND VPWR VPWR _10826_/X sky130_fd_sc_hd__clkbuf_1
X_14594_ _11316_/X _14594_/D VGND VGND VPWR VPWR _14594_/Q sky130_fd_sc_hd__dfxtp_1
X_10757_ _14738_/Q _10749_/X _10756_/X _10752_/X VGND VGND VPWR VPWR _14738_/D sky130_fd_sc_hd__a22o_1
X_13545_ _13544_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13545_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13476_ _13816_/X _13821_/X _13521_/S VGND VGND VPWR VPWR _13476_/X sky130_fd_sc_hd__mux2_2
X_10688_ _14751_/Q _10682_/X _10684_/X _10687_/X VGND VGND VPWR VPWR _14751_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12427_ _12512_/A VGND VGND VPWR VPWR _12428_/A sky130_fd_sc_hd__clkbuf_2
X_15215_ _08868_/X _15215_/D VGND VGND VPWR VPWR _15215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12358_ _12431_/B _12357_/X _12431_/B _12357_/X VGND VGND VPWR VPWR _12358_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_99_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15146_ _09125_/X _15146_/D VGND VGND VPWR VPWR _15146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11309_ _14597_/Q _11303_/X _11195_/X _11304_/X VGND VGND VPWR VPWR _14597_/D sky130_fd_sc_hd__a22o_1
XFILLER_141_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15077_ _09400_/X _15077_/D VGND VGND VPWR VPWR _15077_/Q sky130_fd_sc_hd__dfxtp_1
X_12289_ _12289_/A VGND VGND VPWR VPWR _12289_/Y sky130_fd_sc_hd__inv_2
X_14028_ _14525_/Q _14493_/Q _14461_/Q _14429_/Q _14060_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14028_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08520_ _08520_/A VGND VGND VPWR VPWR _08520_/X sky130_fd_sc_hd__buf_1
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08451_ _08451_/A VGND VGND VPWR VPWR _08451_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07402_ _07402_/A _13543_/X VGND VGND VPWR VPWR _15588_/D sky130_fd_sc_hd__and2_1
X_08382_ _14330_/Q VGND VGND VPWR VPWR _10697_/A sky130_fd_sc_hd__buf_1
XFILLER_149_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07333_ _07337_/A _07333_/B VGND VGND VPWR VPWR _15602_/D sky130_fd_sc_hd__nor2_1
XFILLER_32_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07264_ _07265_/A _07264_/B VGND VGND VPWR VPWR _15626_/D sky130_fd_sc_hd__nor2_1
XFILLER_136_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09003_ _09023_/A VGND VGND VPWR VPWR _09012_/A sky130_fd_sc_hd__buf_1
XFILLER_117_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07195_ _13116_/X _07194_/Y _07191_/X _07177_/B VGND VGND VPWR VPWR _15662_/D sky130_fd_sc_hd__o211a_1
XFILLER_105_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09905_ _14952_/Q _09898_/X _09672_/X _09899_/X VGND VGND VPWR VPWR _14952_/D sky130_fd_sc_hd__a22o_1
X_09836_ _09836_/A VGND VGND VPWR VPWR _09836_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09767_ _09767_/A VGND VGND VPWR VPWR _09767_/X sky130_fd_sc_hd__buf_1
XFILLER_100_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08718_ _08722_/A VGND VGND VPWR VPWR _08718_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09698_ _09724_/A VGND VGND VPWR VPWR _09709_/A sky130_fd_sc_hd__buf_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08649_ _15271_/Q _08647_/X _08523_/X _08648_/X VGND VGND VPWR VPWR _15271_/D sky130_fd_sc_hd__a22o_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ _11755_/A VGND VGND VPWR VPWR _11725_/A sky130_fd_sc_hd__buf_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10611_ _10615_/A VGND VGND VPWR VPWR _10611_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _11612_/A VGND VGND VPWR VPWR _11591_/X sky130_fd_sc_hd__buf_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _13366_/X _13364_/X _13415_/S VGND VGND VPWR VPWR _13330_/X sky130_fd_sc_hd__mux2_1
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10542_ _10542_/A VGND VGND VPWR VPWR _10547_/A sky130_fd_sc_hd__buf_1
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _13260_/X _12452_/B _15565_/Q VGND VGND VPWR VPWR _13261_/X sky130_fd_sc_hd__mux2_1
X_10473_ _10479_/A VGND VGND VPWR VPWR _10473_/X sky130_fd_sc_hd__clkbuf_1
X_12212_ _15564_/Q VGND VGND VPWR VPWR _12867_/A sky130_fd_sc_hd__buf_1
X_15000_ _09739_/X _15000_/D VGND VGND VPWR VPWR _15000_/Q sky130_fd_sc_hd__dfxtp_1
X_13192_ _12395_/A _12329_/X _15561_/Q VGND VGND VPWR VPWR _13192_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12143_ _12138_/X _12287_/B _12142_/Y VGND VGND VPWR VPWR _12636_/A sky130_fd_sc_hd__a21oi_1
XFILLER_2_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12074_ _12065_/X _12092_/A _12599_/A _12094_/A VGND VGND VPWR VPWR _12075_/B sky130_fd_sc_hd__o22a_1
XFILLER_123_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11025_ _11046_/A VGND VGND VPWR VPWR _11025_/X sky130_fd_sc_hd__buf_1
XFILLER_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12976_ _12036_/A _12978_/B _12963_/X _13420_/X _13421_/X VGND VGND VPWR VPWR _12976_/Y
+ sky130_fd_sc_hd__a311oi_4
X_14715_ _10867_/X _14715_/D VGND VGND VPWR VPWR _14715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11927_ _11987_/A VGND VGND VPWR VPWR _11947_/A sky130_fd_sc_hd__buf_2
X_14646_ _11118_/X _14646_/D VGND VGND VPWR VPWR _14646_/Q sky130_fd_sc_hd__dfxtp_1
X_11858_ _14451_/Q _11856_/X _08016_/A _11857_/X VGND VGND VPWR VPWR _14451_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10809_ _11549_/A VGND VGND VPWR VPWR _10809_/X sky130_fd_sc_hd__buf_1
XANTENNA_19 data_address[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14577_ _11381_/X _14577_/D VGND VGND VPWR VPWR _14577_/Q sky130_fd_sc_hd__dfxtp_1
X_11789_ _14470_/Q _11783_/X _11557_/X _11784_/X VGND VGND VPWR VPWR _14470_/D sky130_fd_sc_hd__a22o_1
XFILLER_41_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13528_ _13986_/X _13991_/X _13648_/S VGND VGND VPWR VPWR _13528_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13459_ _13458_/X rdata[21] _13516_/S VGND VGND VPWR VPWR _13459_/X sky130_fd_sc_hd__mux2_2
XFILLER_127_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15129_ _09194_/X _15129_/D VGND VGND VPWR VPWR _15129_/Q sky130_fd_sc_hd__dfxtp_1
X_07951_ _07951_/A VGND VGND VPWR VPWR _07951_/X sky130_fd_sc_hd__clkbuf_2
X_07882_ _07893_/A VGND VGND VPWR VPWR _07882_/X sky130_fd_sc_hd__buf_1
XFILLER_95_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09621_ _10760_/A VGND VGND VPWR VPWR _10375_/A sky130_fd_sc_hd__buf_1
XFILLER_55_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09552_ _10690_/A VGND VGND VPWR VPWR _10320_/A sky130_fd_sc_hd__buf_1
X_08503_ _14311_/Q VGND VGND VPWR VPWR _10798_/A sky130_fd_sc_hd__buf_1
XFILLER_64_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09483_ _15054_/Q _09475_/X _09245_/X _09476_/X VGND VGND VPWR VPWR _15054_/D sky130_fd_sc_hd__a22o_1
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08434_ _09216_/A VGND VGND VPWR VPWR _08434_/X sky130_fd_sc_hd__buf_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08365_ _08481_/A VGND VGND VPWR VPWR _08405_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07316_ _14377_/Q VGND VGND VPWR VPWR _07513_/B sky130_fd_sc_hd__inv_2
XFILLER_109_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08296_ _09000_/A VGND VGND VPWR VPWR _08583_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_109_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07247_ _07247_/A VGND VGND VPWR VPWR _07274_/A sky130_fd_sc_hd__buf_1
XFILLER_118_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07178_ _07252_/B _07190_/A VGND VGND VPWR VPWR _07179_/B sky130_fd_sc_hd__or2_2
XFILLER_118_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09819_ _14977_/Q _09812_/X _09534_/X _09815_/X VGND VGND VPWR VPWR _14977_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12830_ _12830_/A VGND VGND VPWR VPWR _12830_/X sky130_fd_sc_hd__buf_1
X_12761_ _13313_/X VGND VGND VPWR VPWR _12850_/A sky130_fd_sc_hd__inv_2
XFILLER_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14500_ _11681_/X _14500_/D VGND VGND VPWR VPWR _14500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11712_ _11712_/A VGND VGND VPWR VPWR _11712_/X sky130_fd_sc_hd__clkbuf_1
X_12692_ _12692_/A VGND VGND VPWR VPWR _12692_/X sky130_fd_sc_hd__buf_1
XFILLER_42_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15480_ _15509_/CLK _15480_/D VGND VGND VPWR VPWR wdata[6] sky130_fd_sc_hd__dfxtp_2
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11643_ _11643_/A VGND VGND VPWR VPWR _11643_/X sky130_fd_sc_hd__buf_1
X_14431_ _11922_/X _14431_/D VGND VGND VPWR VPWR _14431_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14362_ _15666_/CLK pc[23] VGND VGND VPWR VPWR _14362_/Q sky130_fd_sc_hd__dfxtp_1
X_11574_ _11574_/A _11574_/B _11574_/C VGND VGND VPWR VPWR _11910_/B sky130_fd_sc_hd__or3_1
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _12873_/Y _12927_/Y _13408_/S VGND VGND VPWR VPWR _13313_/X sky130_fd_sc_hd__mux2_1
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10525_ _10531_/A VGND VGND VPWR VPWR _10525_/X sky130_fd_sc_hd__clkbuf_1
X_14293_ _15604_/CLK _15460_/Q VGND VGND VPWR VPWR _14293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13244_ _13245_/X _12823_/A _13393_/S VGND VGND VPWR VPWR _13244_/X sky130_fd_sc_hd__mux2_2
X_10456_ _10475_/A VGND VGND VPWR VPWR _10456_/X sky130_fd_sc_hd__buf_1
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13175_ _13174_/X _13215_/X _13393_/S VGND VGND VPWR VPWR _13175_/X sky130_fd_sc_hd__mux2_1
X_10387_ _10413_/A VGND VGND VPWR VPWR _10398_/A sky130_fd_sc_hd__buf_1
XFILLER_123_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12126_ _15545_/Q VGND VGND VPWR VPWR _12661_/A sky130_fd_sc_hd__inv_2
XFILLER_2_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12057_ _07637_/B _12040_/X _12048_/Y _12031_/X _12056_/Y VGND VGND VPWR VPWR _12307_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_78_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11008_ _14675_/Q _11006_/X _10751_/X _11007_/X VGND VGND VPWR VPWR _14675_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12959_ _12959_/A _12959_/B _12959_/C _12959_/D VGND VGND VPWR VPWR _12963_/A sky130_fd_sc_hd__or4_4
XFILLER_33_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14629_ _11194_/X _14629_/D VGND VGND VPWR VPWR _14629_/Q sky130_fd_sc_hd__dfxtp_1
X_08150_ _08150_/A VGND VGND VPWR VPWR _08159_/A sky130_fd_sc_hd__buf_1
X_08081_ _15399_/Q _08077_/X _08079_/X _08080_/X VGND VGND VPWR VPWR _15399_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08983_ _08989_/A VGND VGND VPWR VPWR _08983_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07934_ _07934_/A VGND VGND VPWR VPWR _07934_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07865_ _07871_/A _07871_/B VGND VGND VPWR VPWR _07872_/B sky130_fd_sc_hd__or2_1
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ _09634_/A VGND VGND VPWR VPWR _09615_/A sky130_fd_sc_hd__buf_1
XFILLER_56_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07796_ _07838_/A VGND VGND VPWR VPWR _07796_/X sky130_fd_sc_hd__buf_1
X_09535_ _15041_/Q _09525_/X _09534_/X _09530_/X VGND VGND VPWR VPWR _15041_/D sky130_fd_sc_hd__a22o_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09466_ _09475_/A VGND VGND VPWR VPWR _09466_/X sky130_fd_sc_hd__buf_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08417_ _08431_/A VGND VGND VPWR VPWR _08417_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09397_ _15079_/Q _09395_/X _09275_/X _09396_/X VGND VGND VPWR VPWR _15079_/D sky130_fd_sc_hd__a22o_1
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08348_ _08364_/A VGND VGND VPWR VPWR _08370_/A sky130_fd_sc_hd__inv_2
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08279_ _08281_/A VGND VGND VPWR VPWR _08279_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10310_ _10319_/A VGND VGND VPWR VPWR _10310_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11290_ _11290_/A VGND VGND VPWR VPWR _11290_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10241_ _10261_/A VGND VGND VPWR VPWR _10246_/A sky130_fd_sc_hd__buf_1
XFILLER_98_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10172_ _14885_/Q _10166_/X _10059_/X _10167_/X VGND VGND VPWR VPWR _14885_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14980_ _09805_/X _14980_/D VGND VGND VPWR VPWR _14980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13931_ _13927_/X _13928_/X _13929_/X _13930_/X _14401_/Q _13966_/S1 VGND VGND VPWR
+ VPWR _13931_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13862_ _15213_/Q _14541_/Q _14989_/Q _15405_/Q _14399_/Q _14400_/Q VGND VGND VPWR
+ VPWR _13862_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15601_ _15601_/CLK _15601_/D VGND VGND VPWR VPWR _15601_/Q sky130_fd_sc_hd__dfxtp_1
X_12813_ _13291_/X _12782_/X _12821_/A _12811_/X _12812_/X VGND VGND VPWR VPWR _12813_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13793_ _14676_/Q _15252_/Q _14740_/Q _14708_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13793_/X sky130_fd_sc_hd__mux4_2
X_15532_ _15578_/CLK _15532_/D VGND VGND VPWR VPWR _15532_/Q sky130_fd_sc_hd__dfxtp_1
X_12744_ _12428_/X _12721_/Y _12735_/X _12743_/Y VGND VGND VPWR VPWR _12744_/X sky130_fd_sc_hd__a31o_1
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15463_ _15604_/CLK _15463_/D VGND VGND VPWR VPWR _15463_/Q sky130_fd_sc_hd__dfxtp_1
X_12675_ _12675_/A VGND VGND VPWR VPWR _12676_/A sky130_fd_sc_hd__buf_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ _11981_/X _14414_/D VGND VGND VPWR VPWR _14414_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _11628_/A VGND VGND VPWR VPWR _11626_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15394_ _08102_/X _15394_/D VGND VGND VPWR VPWR _15394_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ _15648_/CLK pc[6] VGND VGND VPWR VPWR _14345_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11557_ _11557_/A VGND VGND VPWR VPWR _11557_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10508_ _10510_/A VGND VGND VPWR VPWR _10508_/X sky130_fd_sc_hd__clkbuf_1
X_11488_ _11513_/A VGND VGND VPWR VPWR _11488_/X sky130_fd_sc_hd__buf_1
X_14276_ _14272_/X _14273_/X _14274_/X _14275_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14276_/X sky130_fd_sc_hd__mux4_2
X_13227_ _12635_/X _12138_/X _13418_/S VGND VGND VPWR VPWR _13227_/X sky130_fd_sc_hd__mux2_1
Xrepeater7 ren VGND VGND VPWR VPWR _13058_/S sky130_fd_sc_hd__buf_8
X_10439_ _10451_/A VGND VGND VPWR VPWR _10440_/A sky130_fd_sc_hd__buf_1
X_13158_ _12522_/X _12492_/X _15561_/Q VGND VGND VPWR VPWR _13158_/X sky130_fd_sc_hd__mux2_1
X_12109_ _12109_/A _12284_/B VGND VGND VPWR VPWR _12109_/Y sky130_fd_sc_hd__nor2_1
X_13089_ _12515_/Y _15591_/Q _13090_/S VGND VGND VPWR VPWR _13089_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07650_ _07650_/A VGND VGND VPWR VPWR _07689_/A sky130_fd_sc_hd__buf_1
XFILLER_65_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07581_ _07581_/A _13080_/X VGND VGND VPWR VPWR _15495_/D sky130_fd_sc_hd__and2_1
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09320_ _10270_/A VGND VGND VPWR VPWR _09964_/A sky130_fd_sc_hd__buf_1
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09251_ _09251_/A VGND VGND VPWR VPWR _09276_/A sky130_fd_sc_hd__buf_1
X_08202_ _08211_/A VGND VGND VPWR VPWR _08209_/A sky130_fd_sc_hd__buf_1
X_09182_ _09187_/A VGND VGND VPWR VPWR _09182_/X sky130_fd_sc_hd__clkbuf_1
X_08133_ _08139_/A VGND VGND VPWR VPWR _08133_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08064_ _08064_/A VGND VGND VPWR VPWR _08064_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08966_ _08968_/A VGND VGND VPWR VPWR _08966_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07917_ _11428_/A VGND VGND VPWR VPWR _09700_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_69_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08897_ _08897_/A VGND VGND VPWR VPWR _08970_/A sky130_fd_sc_hd__buf_2
XFILLER_56_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07848_ _07848_/A VGND VGND VPWR VPWR _07848_/X sky130_fd_sc_hd__buf_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07779_ _07779_/A _07779_/B _07779_/C VGND VGND VPWR VPWR _07819_/A sky130_fd_sc_hd__and3_1
X_09518_ _09532_/A VGND VGND VPWR VPWR _09518_/X sky130_fd_sc_hd__clkbuf_1
X_10790_ _10790_/A VGND VGND VPWR VPWR _10821_/A sky130_fd_sc_hd__buf_1
XFILLER_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09449_ _09469_/A VGND VGND VPWR VPWR _09454_/A sky130_fd_sc_hd__buf_2
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12460_ _12745_/A VGND VGND VPWR VPWR _12460_/X sky130_fd_sc_hd__buf_2
XFILLER_12_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11411_ _11413_/A VGND VGND VPWR VPWR _11411_/X sky130_fd_sc_hd__clkbuf_1
X_12391_ _12379_/A _12347_/A _12386_/Y _12437_/A VGND VGND VPWR VPWR _12392_/B sky130_fd_sc_hd__o22a_2
X_14130_ _14963_/Q _15059_/Q _15027_/Q _15091_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14130_/X sky130_fd_sc_hd__mux4_1
X_11342_ _11342_/A VGND VGND VPWR VPWR _11342_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11273_ _11273_/A VGND VGND VPWR VPWR _11273_/X sky130_fd_sc_hd__buf_1
X_14061_ _14057_/X _14058_/X _14059_/X _14060_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14061_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13012_ _14356_/Q VGND VGND VPWR VPWR _13012_/Y sky130_fd_sc_hd__inv_2
X_10224_ _14871_/Q _10217_/X _09981_/X _10218_/X VGND VGND VPWR VPWR _14871_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10155_ _10164_/A VGND VGND VPWR VPWR _10162_/A sky130_fd_sc_hd__buf_1
XFILLER_0_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14963_ _09867_/X _14963_/D VGND VGND VPWR VPWR _14963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10086_ _10106_/A VGND VGND VPWR VPWR _10086_/X sky130_fd_sc_hd__buf_1
X_13914_ _15176_/Q _15144_/Q _14760_/Q _14792_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13914_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14894_ _10141_/X _14894_/D VGND VGND VPWR VPWR _14894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13845_ _15119_/Q _15343_/Q _15311_/Q _15279_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13845_/X sky130_fd_sc_hd__mux4_2
X_13776_ _13772_/X _13773_/X _13774_/X _13775_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13776_/X sky130_fd_sc_hd__mux4_2
X_10988_ _10988_/A VGND VGND VPWR VPWR _10993_/A sky130_fd_sc_hd__buf_1
XFILLER_71_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15515_ _15521_/CLK _15515_/D VGND VGND VPWR VPWR _15515_/Q sky130_fd_sc_hd__dfxtp_1
X_12727_ _12727_/A VGND VGND VPWR VPWR _12727_/X sky130_fd_sc_hd__buf_1
XFILLER_31_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15446_ _15652_/CLK _15446_/D VGND VGND VPWR VPWR data_address[19] sky130_fd_sc_hd__dfxtp_4
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ _12371_/A _12656_/Y _13224_/X _12451_/A _12657_/Y VGND VGND VPWR VPWR _12658_/X
+ sky130_fd_sc_hd__o221a_1
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11609_ _14522_/Q _11603_/X _11471_/X _11604_/X VGND VGND VPWR VPWR _14522_/D sky130_fd_sc_hd__a22o_1
XFILLER_129_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15377_ _08169_/X _15377_/D VGND VGND VPWR VPWR _15377_/Q sky130_fd_sc_hd__dfxtp_1
X_12589_ _12588_/X _12079_/X _12360_/X VGND VGND VPWR VPWR _12589_/Y sky130_fd_sc_hd__o21ai_2
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14328_ _14328_/CLK _14328_/D VGND VGND VPWR VPWR _14328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14259_ _14822_/Q _14854_/Q _14886_/Q _14918_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14259_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08820_ _08846_/A VGND VGND VPWR VPWR _08829_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08751_ _15243_/Q _08742_/X _08499_/X _08744_/X VGND VGND VPWR VPWR _15243_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07702_ _07701_/X _13135_/X _07681_/X VGND VGND VPWR VPWR _07852_/A sky130_fd_sc_hd__a21bo_1
X_08682_ _08703_/A VGND VGND VPWR VPWR _08682_/X sky130_fd_sc_hd__buf_1
XFILLER_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07633_ _07634_/A _07633_/B VGND VGND VPWR VPWR _15466_/D sky130_fd_sc_hd__nor2_1
XFILLER_81_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07564_ _13648_/S _07530_/Y _14398_/Q _07540_/Y _07563_/X VGND VGND VPWR VPWR _07564_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09303_ _09305_/A VGND VGND VPWR VPWR _09303_/X sky130_fd_sc_hd__clkbuf_1
X_07495_ _07495_/A _07495_/B VGND VGND VPWR VPWR _15524_/D sky130_fd_sc_hd__nor2_1
XFILLER_139_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09234_ _09239_/A VGND VGND VPWR VPWR _09234_/X sky130_fd_sc_hd__clkbuf_1
X_09165_ _15136_/Q _09152_/X _09164_/X _09156_/X VGND VGND VPWR VPWR _15136_/D sky130_fd_sc_hd__a22o_1
X_08116_ _08116_/A VGND VGND VPWR VPWR _08116_/X sky130_fd_sc_hd__clkbuf_1
X_09096_ _09107_/A VGND VGND VPWR VPWR _09096_/X sky130_fd_sc_hd__buf_1
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08047_ _14314_/Q VGND VGND VPWR VPWR _08048_/A sky130_fd_sc_hd__buf_1
XFILLER_89_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09998_ _10011_/A VGND VGND VPWR VPWR _09998_/X sky130_fd_sc_hd__buf_1
XFILLER_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08949_ _15198_/Q _08943_/X _08805_/X _08946_/X VGND VGND VPWR VPWR _15198_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11960_ _11962_/A VGND VGND VPWR VPWR _11960_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10911_ _10922_/A VGND VGND VPWR VPWR _10920_/A sky130_fd_sc_hd__buf_1
XFILLER_45_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11891_ _11900_/A VGND VGND VPWR VPWR _11898_/A sky130_fd_sc_hd__buf_1
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13630_ _13629_/X _14309_/D _15506_/Q VGND VGND VPWR VPWR _13630_/X sky130_fd_sc_hd__mux2_1
X_10842_ _10854_/A VGND VGND VPWR VPWR _10843_/A sky130_fd_sc_hd__buf_1
XFILLER_60_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13561_ _13560_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13561_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10773_ _10773_/A VGND VGND VPWR VPWR _10786_/A sky130_fd_sc_hd__buf_2
X_15300_ _08537_/X _15300_/D VGND VGND VPWR VPWR _15300_/Q sky130_fd_sc_hd__dfxtp_1
X_12512_ _12512_/A VGND VGND VPWR VPWR _12512_/X sky130_fd_sc_hd__clkbuf_4
X_13492_ _13491_/X rdata[10] _13516_/S VGND VGND VPWR VPWR _13492_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15231_ _08795_/X _15231_/D VGND VGND VPWR VPWR _15231_/Q sky130_fd_sc_hd__dfxtp_1
X_12443_ _12443_/A _12443_/B VGND VGND VPWR VPWR _12443_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15162_ _09072_/X _15162_/D VGND VGND VPWR VPWR _15162_/Q sky130_fd_sc_hd__dfxtp_1
X_12374_ _12368_/X _12345_/X _12371_/X _12373_/Y VGND VGND VPWR VPWR _12374_/X sky130_fd_sc_hd__o22a_1
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14113_ _14676_/Q _15252_/Q _14740_/Q _14708_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14113_/X sky130_fd_sc_hd__mux4_2
X_11325_ _11329_/A VGND VGND VPWR VPWR _11325_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15093_ _09349_/X _15093_/D VGND VGND VPWR VPWR _15093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14044_ _15195_/Q _15163_/Q _14779_/Q _14811_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14044_/X sky130_fd_sc_hd__mux4_2
X_11256_ _11274_/A VGND VGND VPWR VPWR _11256_/X sky130_fd_sc_hd__buf_1
XFILLER_69_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10207_ _10217_/A VGND VGND VPWR VPWR _10207_/X sky130_fd_sc_hd__buf_1
X_11187_ _11553_/A VGND VGND VPWR VPWR _11187_/X sky130_fd_sc_hd__buf_1
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10138_ _14896_/Q _10136_/X _10012_/X _10137_/X VGND VGND VPWR VPWR _14896_/D sky130_fd_sc_hd__a22o_1
XFILLER_94_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10069_ _10548_/A _10181_/B VGND VGND VPWR VPWR _10084_/A sky130_fd_sc_hd__or2_2
X_14946_ _09921_/X _14946_/D VGND VGND VPWR VPWR _14946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14877_ _10204_/X _14877_/D VGND VGND VPWR VPWR _14877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13828_ _14513_/Q _14481_/Q _14449_/Q _14417_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13828_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13759_ _14840_/Q _14872_/Q _14904_/Q _14936_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13759_/X sky130_fd_sc_hd__mux4_2
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07280_ _07282_/A _07280_/B VGND VGND VPWR VPWR _15615_/D sky130_fd_sc_hd__nor2_1
XFILLER_148_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15429_ _15604_/CLK _15429_/D VGND VGND VPWR VPWR data_address[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_116_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09921_ _09933_/A VGND VGND VPWR VPWR _09921_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09852_ _09854_/A VGND VGND VPWR VPWR _09852_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08803_ _15231_/Q _08798_/X _08799_/X _08802_/X VGND VGND VPWR VPWR _15231_/D sky130_fd_sc_hd__a22o_1
X_09783_ _09783_/A VGND VGND VPWR VPWR _09783_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08734_ _15248_/Q _08732_/X _08466_/X _08733_/X VGND VGND VPWR VPWR _15248_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_109 pc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08665_ _08677_/A VGND VGND VPWR VPWR _08666_/A sky130_fd_sc_hd__buf_1
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07616_ _12049_/A VGND VGND VPWR VPWR _07617_/A sky130_fd_sc_hd__inv_2
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08596_ _08626_/A VGND VGND VPWR VPWR _08617_/A sky130_fd_sc_hd__clkbuf_2
X_07547_ _15514_/Q VGND VGND VPWR VPWR _07633_/B sky130_fd_sc_hd__inv_2
XFILLER_10_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07478_ _07478_/A _13499_/X VGND VGND VPWR VPWR _15537_/D sky130_fd_sc_hd__and2_1
XFILLER_22_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09217_ _15125_/Q _09210_/X _09216_/X _09213_/X VGND VGND VPWR VPWR _15125_/D sky130_fd_sc_hd__a22o_1
X_09148_ _15139_/Q _09041_/A _08919_/X _09044_/A VGND VGND VPWR VPWR _15139_/D sky130_fd_sc_hd__a22o_1
XFILLER_107_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09079_ _09083_/A VGND VGND VPWR VPWR _09079_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11110_ _14649_/Q _11107_/X _11108_/X _11109_/X VGND VGND VPWR VPWR _14649_/D sky130_fd_sc_hd__a22o_1
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12090_ _15549_/Q VGND VGND VPWR VPWR _12611_/A sky130_fd_sc_hd__inv_2
X_11041_ _11045_/A VGND VGND VPWR VPWR _11041_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14800_ _10504_/X _14800_/D VGND VGND VPWR VPWR _14800_/Q sky130_fd_sc_hd__dfxtp_1
X_12992_ _12988_/X _12991_/X _12993_/B VGND VGND VPWR VPWR _12992_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14731_ _10792_/X _14731_/D VGND VGND VPWR VPWR _14731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11943_ _11973_/A VGND VGND VPWR VPWR _11964_/A sky130_fd_sc_hd__buf_2
XFILLER_72_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14662_ _11050_/X _14662_/D VGND VGND VPWR VPWR _14662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11874_ _11874_/A VGND VGND VPWR VPWR _11895_/A sky130_fd_sc_hd__clkbuf_2
X_13613_ _13612_/X _07332_/Y _13649_/S VGND VGND VPWR VPWR _13613_/X sky130_fd_sc_hd__mux2_1
X_10825_ _14725_/Q _10812_/X _10824_/X _10815_/X VGND VGND VPWR VPWR _14725_/D sky130_fd_sc_hd__a22o_1
X_14593_ _11325_/X _14593_/D VGND VGND VPWR VPWR _14593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13544_ _14026_/X _14031_/X _14387_/Q VGND VGND VPWR VPWR _13544_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10756_ _11506_/A VGND VGND VPWR VPWR _10756_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13475_ _13474_/X _13075_/X _14336_/Q VGND VGND VPWR VPWR _13475_/X sky130_fd_sc_hd__mux2_1
X_10687_ _10719_/A VGND VGND VPWR VPWR _10687_/X sky130_fd_sc_hd__buf_1
XFILLER_145_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15214_ _08872_/X _15214_/D VGND VGND VPWR VPWR _15214_/Q sky130_fd_sc_hd__dfxtp_1
X_12426_ _12426_/A VGND VGND VPWR VPWR _12512_/A sky130_fd_sc_hd__inv_2
XFILLER_65_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15145_ _09131_/X _15145_/D VGND VGND VPWR VPWR _15145_/Q sky130_fd_sc_hd__dfxtp_1
X_12357_ _12357_/A _12357_/B VGND VGND VPWR VPWR _12357_/X sky130_fd_sc_hd__or2_1
XFILLER_5_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11308_ _11308_/A VGND VGND VPWR VPWR _11308_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15076_ _09403_/X _15076_/D VGND VGND VPWR VPWR _15076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12288_ _15545_/Q _12133_/Y _12287_/Y _12142_/Y VGND VGND VPWR VPWR _12289_/A sky130_fd_sc_hd__a31o_1
X_14027_ _14653_/Q _14621_/Q _14589_/Q _15389_/Q _14060_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14027_/X sky130_fd_sc_hd__mux4_2
XFILLER_68_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11239_ _11239_/A VGND VGND VPWR VPWR _11246_/A sky130_fd_sc_hd__buf_1
XFILLER_122_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14929_ _10007_/X _14929_/D VGND VGND VPWR VPWR _14929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08450_ _15315_/Q _08445_/X _08448_/X _08449_/X VGND VGND VPWR VPWR _15315_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07401_ _07402_/A _13539_/X VGND VGND VPWR VPWR _15589_/D sky130_fd_sc_hd__and2_1
X_08381_ _08393_/A VGND VGND VPWR VPWR _08381_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07332_ _07333_/B VGND VGND VPWR VPWR _07332_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07263_ _07265_/A _07263_/B VGND VGND VPWR VPWR _15627_/D sky130_fd_sc_hd__nor2_1
XFILLER_118_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09002_ _09068_/A VGND VGND VPWR VPWR _09023_/A sky130_fd_sc_hd__clkbuf_2
X_07194_ _07194_/A VGND VGND VPWR VPWR _07194_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09904_ _09906_/A VGND VGND VPWR VPWR _09904_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09835_ _14973_/Q _09825_/X _09559_/X _09828_/X VGND VGND VPWR VPWR _14973_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09766_ _09772_/A VGND VGND VPWR VPWR _09766_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08717_ _08735_/A VGND VGND VPWR VPWR _08722_/A sky130_fd_sc_hd__buf_1
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09697_ _09733_/A VGND VGND VPWR VPWR _09724_/A sky130_fd_sc_hd__clkbuf_4
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08648_ _08648_/A VGND VGND VPWR VPWR _08648_/X sky130_fd_sc_hd__buf_1
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08579_ _08581_/A VGND VGND VPWR VPWR _08579_/X sky130_fd_sc_hd__clkbuf_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10610_ _10610_/A VGND VGND VPWR VPWR _10615_/A sky130_fd_sc_hd__buf_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11590_ _11651_/A VGND VGND VPWR VPWR _11612_/A sky130_fd_sc_hd__buf_2
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ _14789_/Q _10535_/X _10428_/X _10536_/X VGND VGND VPWR VPWR _14789_/D sky130_fd_sc_hd__a22o_1
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13260_ _13321_/X _13320_/X _13393_/S VGND VGND VPWR VPWR _13260_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10472_ _10481_/A VGND VGND VPWR VPWR _10479_/A sky130_fd_sc_hd__buf_1
X_12211_ _12230_/A VGND VGND VPWR VPWR _12211_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13191_ _13192_/X _13202_/X _15562_/Q VGND VGND VPWR VPWR _13191_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12142_ _12142_/A _12287_/B VGND VGND VPWR VPWR _12142_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12073_ _12105_/A VGND VGND VPWR VPWR _12094_/A sky130_fd_sc_hd__buf_1
XFILLER_123_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11024_ _11024_/A VGND VGND VPWR VPWR _11046_/A sky130_fd_sc_hd__buf_1
XFILLER_37_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12975_ _12975_/A VGND VGND VPWR VPWR _12978_/B sky130_fd_sc_hd__inv_2
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14714_ _10869_/X _14714_/D VGND VGND VPWR VPWR _14714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11926_ _11926_/A VGND VGND VPWR VPWR _11987_/A sky130_fd_sc_hd__buf_2
XFILLER_18_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14645_ _11125_/X _14645_/D VGND VGND VPWR VPWR _14645_/Q sky130_fd_sc_hd__dfxtp_1
X_11857_ _11866_/A VGND VGND VPWR VPWR _11857_/X sky130_fd_sc_hd__buf_1
XFILLER_82_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10808_ _10808_/A VGND VGND VPWR VPWR _11549_/A sky130_fd_sc_hd__clkbuf_2
X_14576_ _11383_/X _14576_/D VGND VGND VPWR VPWR _14576_/Q sky130_fd_sc_hd__dfxtp_1
X_11788_ _11792_/A VGND VGND VPWR VPWR _11788_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13527_ _13526_/X _13090_/X _14337_/Q VGND VGND VPWR VPWR _13527_/X sky130_fd_sc_hd__mux2_1
X_10739_ _10739_/A VGND VGND VPWR VPWR _11494_/A sky130_fd_sc_hd__clkbuf_2
X_13458_ _13756_/X _13761_/X _13521_/S VGND VGND VPWR VPWR _13458_/X sky130_fd_sc_hd__mux2_1
X_12409_ _12409_/A VGND VGND VPWR VPWR _12432_/B sky130_fd_sc_hd__inv_2
X_13389_ _13388_/X _13418_/X _13415_/S VGND VGND VPWR VPWR _13389_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15128_ _09199_/X _15128_/D VGND VGND VPWR VPWR _15128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15059_ _09465_/X _15059_/D VGND VGND VPWR VPWR _15059_/Q sky130_fd_sc_hd__dfxtp_1
X_07950_ _14332_/Q VGND VGND VPWR VPWR _07951_/A sky130_fd_sc_hd__buf_1
XFILLER_102_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07881_ _07772_/A _07880_/Y _07722_/A _07880_/A _07869_/X VGND VGND VPWR VPWR _15438_/D
+ sky130_fd_sc_hd__o221a_1
X_09620_ _09630_/A VGND VGND VPWR VPWR _09620_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09551_ _09551_/A VGND VGND VPWR VPWR _09551_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08502_ _08520_/A VGND VGND VPWR VPWR _08502_/X sky130_fd_sc_hd__buf_1
XFILLER_24_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09482_ _09484_/A VGND VGND VPWR VPWR _09482_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08433_ _10739_/A VGND VGND VPWR VPWR _09216_/A sky130_fd_sc_hd__buf_1
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08364_ _08364_/A VGND VGND VPWR VPWR _08481_/A sky130_fd_sc_hd__buf_4
X_07315_ _14378_/Q VGND VGND VPWR VPWR _07512_/B sky130_fd_sc_hd__inv_2
X_08295_ _10270_/A VGND VGND VPWR VPWR _09000_/A sky130_fd_sc_hd__buf_1
XFILLER_20_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07246_ _07246_/A _07246_/B VGND VGND VPWR VPWR _15637_/D sky130_fd_sc_hd__or2_1
X_07177_ _07254_/B _07177_/B VGND VGND VPWR VPWR _07190_/A sky130_fd_sc_hd__or2_1
XFILLER_133_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09818_ _09822_/A VGND VGND VPWR VPWR _09818_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09749_ _14998_/Q _09746_/X _09595_/X _09748_/X VGND VGND VPWR VPWR _14998_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12760_ _12745_/X _12751_/Y _12757_/Y _12759_/X VGND VGND VPWR VPWR _12760_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_55_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11711_ _14493_/Q _11702_/X _11459_/X _11705_/X VGND VGND VPWR VPWR _14493_/D sky130_fd_sc_hd__a22o_1
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12162_/A _12690_/X _12162_/A _12690_/X VGND VGND VPWR VPWR _12691_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_70_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _11930_/X _14430_/D VGND VGND VPWR VPWR _14430_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11642_/A VGND VGND VPWR VPWR _11642_/X sky130_fd_sc_hd__buf_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _15621_/CLK pc[22] VGND VGND VPWR VPWR _14361_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11573_ _11585_/A VGND VGND VPWR VPWR _11573_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _13376_/X _13372_/X _13408_/S VGND VGND VPWR VPWR _13312_/X sky130_fd_sc_hd__mux2_1
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10524_ _10542_/A VGND VGND VPWR VPWR _10531_/A sky130_fd_sc_hd__buf_1
X_14292_ _15604_/CLK _15459_/Q VGND VGND VPWR VPWR _14292_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13243_ _13242_/X _12521_/X _15565_/Q VGND VGND VPWR VPWR _13243_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10455_ _10516_/A VGND VGND VPWR VPWR _10475_/A sky130_fd_sc_hd__clkbuf_2
X_13174_ _13173_/X _13196_/X _13408_/S VGND VGND VPWR VPWR _13174_/X sky130_fd_sc_hd__mux2_1
X_10386_ _10462_/A VGND VGND VPWR VPWR _10413_/A sky130_fd_sc_hd__buf_1
XFILLER_97_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12125_ _12640_/A _12651_/A VGND VGND VPWR VPWR _12144_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12056_ _13425_/S _12055_/Y _12024_/X VGND VGND VPWR VPWR _12056_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11007_ _11016_/A VGND VGND VPWR VPWR _11007_/X sky130_fd_sc_hd__buf_1
XFILLER_78_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12958_ _12958_/A _12958_/B VGND VGND VPWR VPWR _12959_/B sky130_fd_sc_hd__or2_1
XFILLER_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11909_ _11919_/A VGND VGND VPWR VPWR _11909_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12889_ _12886_/X _12885_/X _12830_/X VGND VGND VPWR VPWR _12889_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14628_ _11197_/X _14628_/D VGND VGND VPWR VPWR _14628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14559_ _11445_/X _14559_/D VGND VGND VPWR VPWR _14559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08080_ _08080_/A VGND VGND VPWR VPWR _08080_/X sky130_fd_sc_hd__buf_1
XFILLER_146_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08982_ _08991_/A VGND VGND VPWR VPWR _08989_/A sky130_fd_sc_hd__buf_1
XFILLER_114_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07933_ _15426_/Q _07927_/X _07929_/X _07932_/X VGND VGND VPWR VPWR _15426_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07864_ _07872_/A _07864_/B _07864_/C VGND VGND VPWR VPWR _15441_/D sky130_fd_sc_hd__and3_1
XFILLER_95_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09603_ _09603_/A VGND VGND VPWR VPWR _09634_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07795_ _07795_/A VGND VGND VPWR VPWR _07838_/A sky130_fd_sc_hd__buf_1
XFILLER_37_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09534_ _10303_/A VGND VGND VPWR VPWR _09534_/X sky130_fd_sc_hd__buf_1
XFILLER_43_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09465_ _09465_/A VGND VGND VPWR VPWR _09465_/X sky130_fd_sc_hd__clkbuf_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08416_ _08416_/A VGND VGND VPWR VPWR _08431_/A sky130_fd_sc_hd__clkbuf_4
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09396_ _09396_/A VGND VGND VPWR VPWR _09396_/X sky130_fd_sc_hd__buf_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08347_ _09153_/A VGND VGND VPWR VPWR _08347_/X sky130_fd_sc_hd__buf_1
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08278_ _15349_/Q _08272_/X _08006_/X _08274_/X VGND VGND VPWR VPWR _15349_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07229_ _13098_/X _07228_/Y _07221_/X _07159_/B VGND VGND VPWR VPWR _15644_/D sky130_fd_sc_hd__o211a_1
XFILLER_152_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10240_ _10240_/A VGND VGND VPWR VPWR _10261_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_133_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10171_ _10171_/A VGND VGND VPWR VPWR _10171_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13930_ _14951_/Q _15047_/Q _15015_/Q _15079_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13930_/X sky130_fd_sc_hd__mux4_2
XFILLER_47_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13861_ _13857_/X _13858_/X _13859_/X _13860_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13861_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15600_ _15601_/CLK _15600_/D VGND VGND VPWR VPWR _15600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12812_ _12812_/A _12812_/B _12847_/C VGND VGND VPWR VPWR _12812_/X sky130_fd_sc_hd__or3_1
X_13792_ _15220_/Q _14548_/Q _14996_/Q _15412_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13792_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15531_ _15578_/CLK _15531_/D VGND VGND VPWR VPWR _15531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12743_ _13256_/X _12707_/A _12913_/A _12738_/X _12742_/X VGND VGND VPWR VPWR _12743_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_70_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15462_ _15510_/CLK _15462_/D VGND VGND VPWR VPWR _15462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12663_/X _12665_/Y _12667_/Y _12669_/X _12673_/X VGND VGND VPWR VPWR _12674_/Y
+ sky130_fd_sc_hd__o2111ai_4
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _11984_/X _14413_/D VGND VGND VPWR VPWR _14413_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _14518_/Q _11622_/X _11489_/X _11624_/X VGND VGND VPWR VPWR _14518_/D sky130_fd_sc_hd__a22o_1
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _08114_/X _15393_/D VGND VGND VPWR VPWR _15393_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14344_ _15669_/CLK pc[5] VGND VGND VPWR VPWR _14344_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _11556_/A VGND VGND VPWR VPWR _11556_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10507_ _14800_/Q _10505_/X _10379_/X _10506_/X VGND VGND VPWR VPWR _14800_/D sky130_fd_sc_hd__a22o_1
X_14275_ _15108_/Q _15332_/Q _15300_/Q _15268_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14275_/X sky130_fd_sc_hd__mux4_1
X_11487_ _11526_/A VGND VGND VPWR VPWR _11513_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13226_ _13227_/X _13237_/X _13415_/S VGND VGND VPWR VPWR _13226_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater8 _15564_/Q VGND VGND VPWR VPWR _13393_/S sky130_fd_sc_hd__clkbuf_16
X_10438_ _10838_/A _10438_/B VGND VGND VPWR VPWR _10451_/A sky130_fd_sc_hd__or2_2
XFILLER_124_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13157_ _12568_/Y _07387_/A _13157_/S VGND VGND VPWR VPWR _13157_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10369_ _14835_/Q _10366_/X _10367_/X _10368_/X VGND VGND VPWR VPWR _14835_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12108_ _12101_/X _12346_/A _12618_/A _12300_/A VGND VGND VPWR VPWR _12284_/B sky130_fd_sc_hd__o22a_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13088_ _12482_/Y _15590_/Q _13090_/S VGND VGND VPWR VPWR _13088_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12039_ _15523_/Q _15522_/Q _12039_/C VGND VGND VPWR VPWR _12983_/C sky130_fd_sc_hd__or3_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07580_ _07581_/A _13081_/X VGND VGND VPWR VPWR _15496_/D sky130_fd_sc_hd__and2_1
XFILLER_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09250_ _09250_/A VGND VGND VPWR VPWR _09250_/X sky130_fd_sc_hd__buf_1
XFILLER_33_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08201_ _15368_/Q _08195_/X _08074_/X _08196_/X VGND VGND VPWR VPWR _15368_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09181_ _15133_/Q _09169_/X _09180_/X _09173_/X VGND VGND VPWR VPWR _15133_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08132_ _08150_/A VGND VGND VPWR VPWR _08139_/A sky130_fd_sc_hd__buf_1
XFILLER_147_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08063_ _14311_/Q VGND VGND VPWR VPWR _08064_/A sky130_fd_sc_hd__buf_1
XFILLER_147_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08965_ _15193_/Q _08963_/X _08826_/X _08964_/X VGND VGND VPWR VPWR _15193_/D sky130_fd_sc_hd__a22o_1
XFILLER_76_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07916_ _08925_/A _11574_/B _08925_/C VGND VGND VPWR VPWR _11428_/A sky130_fd_sc_hd__or3_1
X_08896_ _15209_/Q _08890_/X _08895_/X _08892_/X VGND VGND VPWR VPWR _15209_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07847_ _07777_/C _07846_/Y _07838_/X _07841_/X VGND VGND VPWR VPWR _15445_/D sky130_fd_sc_hd__o211a_1
XFILLER_83_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07778_ _07830_/A _07827_/A _07778_/C _07821_/A VGND VGND VPWR VPWR _07779_/C sky130_fd_sc_hd__or4b_1
XFILLER_37_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09517_ _09536_/A VGND VGND VPWR VPWR _09532_/A sky130_fd_sc_hd__buf_1
XFILLER_71_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _09478_/A VGND VGND VPWR VPWR _09469_/A sky130_fd_sc_hd__buf_2
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09379_ _09381_/A VGND VGND VPWR VPWR _09379_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11410_ _14569_/Q _11404_/X _11178_/X _11405_/X VGND VGND VPWR VPWR _14569_/D sky130_fd_sc_hd__a22o_1
X_12390_ _12386_/Y _12388_/X _12365_/X _12389_/X _12376_/X VGND VGND VPWR VPWR _12390_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11341_ _14589_/Q _11332_/X _11091_/X _11335_/X VGND VGND VPWR VPWR _14589_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14060_ _14970_/Q _15066_/Q _15034_/Q _15098_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _14060_/X sky130_fd_sc_hd__mux4_2
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11272_ _11278_/A VGND VGND VPWR VPWR _11272_/X sky130_fd_sc_hd__clkbuf_1
X_13011_ _14355_/Q VGND VGND VPWR VPWR _13011_/Y sky130_fd_sc_hd__inv_2
X_10223_ _10225_/A VGND VGND VPWR VPWR _10223_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10154_ _14891_/Q _10147_/X _10034_/X _10149_/X VGND VGND VPWR VPWR _14891_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14962_ _09872_/X _14962_/D VGND VGND VPWR VPWR _14962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10085_ _10146_/A VGND VGND VPWR VPWR _10106_/A sky130_fd_sc_hd__buf_2
XFILLER_59_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13913_ _14664_/Q _15240_/Q _14728_/Q _14696_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13913_/X sky130_fd_sc_hd__mux4_2
X_14893_ _10145_/X _14893_/D VGND VGND VPWR VPWR _14893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13844_ _15183_/Q _15151_/Q _14767_/Q _14799_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13844_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13775_ _15126_/Q _15350_/Q _15318_/Q _15286_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13775_/X sky130_fd_sc_hd__mux4_1
X_10987_ _14681_/Q _10985_/X _10718_/X _10986_/X VGND VGND VPWR VPWR _14681_/D sky130_fd_sc_hd__a22o_1
XFILLER_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12726_ _12726_/A VGND VGND VPWR VPWR _12730_/B sky130_fd_sc_hd__buf_1
X_15514_ _15527_/CLK _15514_/D VGND VGND VPWR VPWR _15514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15445_ _15654_/CLK _15445_/D VGND VGND VPWR VPWR data_address[18] sky130_fd_sc_hd__dfxtp_4
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ _12120_/X _12654_/X _12829_/A VGND VGND VPWR VPWR _12657_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ _11608_/A VGND VGND VPWR VPWR _11608_/X sky130_fd_sc_hd__clkbuf_1
X_15376_ _08172_/X _15376_/D VGND VGND VPWR VPWR _15376_/Q sky130_fd_sc_hd__dfxtp_1
X_12588_ _12588_/A VGND VGND VPWR VPWR _12588_/X sky130_fd_sc_hd__buf_1
XFILLER_128_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14327_ _15498_/CLK _14327_/D VGND VGND VPWR VPWR _14327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11539_ _11544_/A VGND VGND VPWR VPWR _11539_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14258_ _14502_/Q _14470_/Q _14438_/Q _14406_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14258_/X sky130_fd_sc_hd__mux4_2
XFILLER_143_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13209_ _13208_/X _12846_/X _15565_/Q VGND VGND VPWR VPWR _13209_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14189_ _14829_/Q _14861_/Q _14893_/Q _14925_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14189_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08750_ _08752_/A VGND VGND VPWR VPWR _08750_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07701_ _07701_/A VGND VGND VPWR VPWR _07701_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08681_ _08743_/A VGND VGND VPWR VPWR _08703_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07632_ _07634_/A _07632_/B VGND VGND VPWR VPWR _15467_/D sky130_fd_sc_hd__nor2_1
XFILLER_38_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07563_ _12574_/A _15470_/Q _12569_/A _15467_/Q VGND VGND VPWR VPWR _07563_/X sky130_fd_sc_hd__o22a_1
X_09302_ _15106_/Q _09298_/X _09153_/X _09301_/X VGND VGND VPWR VPWR _15106_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07494_ _07495_/A _07494_/B VGND VGND VPWR VPWR _15525_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09233_ _15121_/Q _09223_/X _09232_/X _09225_/X VGND VGND VPWR VPWR _15121_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09164_ _09164_/A VGND VGND VPWR VPWR _09164_/X sky130_fd_sc_hd__buf_1
XFILLER_108_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08115_ _15393_/Q _08109_/X _07936_/X _08112_/X VGND VGND VPWR VPWR _15393_/D sky130_fd_sc_hd__a22o_1
X_09095_ _09106_/A VGND VGND VPWR VPWR _09095_/X sky130_fd_sc_hd__buf_1
XFILLER_108_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08046_ _08077_/A VGND VGND VPWR VPWR _08046_/X sky130_fd_sc_hd__buf_1
XFILLER_103_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09997_ _10002_/A VGND VGND VPWR VPWR _09997_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08948_ _08950_/A VGND VGND VPWR VPWR _08948_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08879_ _08879_/A VGND VGND VPWR VPWR _08906_/A sky130_fd_sc_hd__buf_1
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10910_ _14702_/Q _10904_/X _10776_/X _10905_/X VGND VGND VPWR VPWR _14702_/D sky130_fd_sc_hd__a22o_1
X_11890_ _14441_/Q _11886_/X _08069_/A _11887_/X VGND VGND VPWR VPWR _14441_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10841_ _10851_/A VGND VGND VPWR VPWR _10854_/A sky130_fd_sc_hd__inv_2
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13560_ _14066_/X _14071_/X _13648_/S VGND VGND VPWR VPWR _13560_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10772_ _14735_/Q _10764_/X _10771_/X _10767_/X VGND VGND VPWR VPWR _14735_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12511_ _12443_/B _12467_/Y _12443_/A _12510_/X VGND VGND VPWR VPWR _12513_/B sky130_fd_sc_hd__a31o_1
X_13491_ _13866_/X _13871_/X _13521_/S VGND VGND VPWR VPWR _13491_/X sky130_fd_sc_hd__mux2_4
XFILLER_8_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15230_ _08804_/X _15230_/D VGND VGND VPWR VPWR _15230_/Q sky130_fd_sc_hd__dfxtp_1
X_12442_ _12443_/A _12443_/B VGND VGND VPWR VPWR _12442_/X sky130_fd_sc_hd__or2_1
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15161_ _09074_/X _15161_/D VGND VGND VPWR VPWR _15161_/Q sky130_fd_sc_hd__dfxtp_1
X_12373_ _12904_/C VGND VGND VPWR VPWR _12373_/Y sky130_fd_sc_hd__inv_2
X_14112_ _15220_/Q _14548_/Q _14996_/Q _15412_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14112_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11324_ _11337_/A VGND VGND VPWR VPWR _11329_/A sky130_fd_sc_hd__buf_1
X_15092_ _09351_/X _15092_/D VGND VGND VPWR VPWR _15092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14043_ _14683_/Q _15259_/Q _14747_/Q _14715_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14043_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11255_ _11285_/A VGND VGND VPWR VPWR _11274_/A sky130_fd_sc_hd__buf_2
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10206_ _10206_/A VGND VGND VPWR VPWR _10206_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11186_ _11186_/A VGND VGND VPWR VPWR _11186_/X sky130_fd_sc_hd__buf_1
XFILLER_122_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10137_ _10137_/A VGND VGND VPWR VPWR _10137_/X sky130_fd_sc_hd__buf_1
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10068_ _10078_/A VGND VGND VPWR VPWR _10068_/X sky130_fd_sc_hd__clkbuf_1
X_14945_ _09933_/X _14945_/D VGND VGND VPWR VPWR _14945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14876_ _10206_/X _14876_/D VGND VGND VPWR VPWR _14876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13827_ _14641_/Q _14609_/Q _14577_/Q _15377_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13827_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13758_ _14520_/Q _14488_/Q _14456_/Q _14424_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13758_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12709_ _12709_/A VGND VGND VPWR VPWR _12709_/X sky130_fd_sc_hd__buf_2
XFILLER_148_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13689_ _14847_/Q _14879_/Q _14911_/Q _14943_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13689_/X sky130_fd_sc_hd__mux4_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15428_ _15601_/CLK _15428_/D VGND VGND VPWR VPWR data_address[1] sky130_fd_sc_hd__dfxtp_2
X_15359_ _08238_/X _15359_/D VGND VGND VPWR VPWR _15359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09920_ _14947_/Q _09812_/A _09695_/X _09815_/A VGND VGND VPWR VPWR _14947_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09851_ _14968_/Q _09846_/X _09584_/X _09847_/X VGND VGND VPWR VPWR _14968_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08802_ _08827_/A VGND VGND VPWR VPWR _08802_/X sky130_fd_sc_hd__buf_1
XFILLER_58_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09782_ _14988_/Q _09777_/X _09649_/X _09779_/X VGND VGND VPWR VPWR _14988_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08733_ _08733_/A VGND VGND VPWR VPWR _08733_/X sky130_fd_sc_hd__buf_1
XFILLER_82_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08664_ _09408_/A _10949_/A VGND VGND VPWR VPWR _08677_/A sky130_fd_sc_hd__or2_2
XFILLER_54_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07615_ _15521_/Q VGND VGND VPWR VPWR _12049_/A sky130_fd_sc_hd__buf_1
XFILLER_81_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08595_ _08603_/A VGND VGND VPWR VPWR _08595_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07546_ _15518_/Q VGND VGND VPWR VPWR _07628_/B sky130_fd_sc_hd__inv_2
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07477_ _07478_/A _13496_/X VGND VGND VPWR VPWR _15538_/D sky130_fd_sc_hd__and2_1
XFILLER_139_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09216_ _09216_/A VGND VGND VPWR VPWR _09216_/X sky130_fd_sc_hd__buf_1
XFILLER_148_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09147_ _09158_/A VGND VGND VPWR VPWR _09147_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09078_ _09089_/A VGND VGND VPWR VPWR _09083_/A sky130_fd_sc_hd__buf_2
XFILLER_108_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08029_ _08029_/A VGND VGND VPWR VPWR _08029_/X sky130_fd_sc_hd__buf_1
XFILLER_150_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11040_ _11049_/A VGND VGND VPWR VPWR _11045_/A sky130_fd_sc_hd__buf_1
XFILLER_122_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12991_ _15515_/Q _12570_/A _07629_/B _14398_/Q _12990_/X VGND VGND VPWR VPWR _12991_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14730_ _10796_/X _14730_/D VGND VGND VPWR VPWR _14730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11942_ _14426_/Q _11936_/X _07978_/A _11937_/X VGND VGND VPWR VPWR _14426_/D sky130_fd_sc_hd__a22o_1
X_14661_ _11052_/X _14661_/D VGND VGND VPWR VPWR _14661_/Q sky130_fd_sc_hd__dfxtp_1
X_11873_ _11879_/A VGND VGND VPWR VPWR _11873_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13612_ _14196_/X _14201_/X _13648_/S VGND VGND VPWR VPWR _13612_/X sky130_fd_sc_hd__mux2_4
X_10824_ _11564_/A VGND VGND VPWR VPWR _10824_/X sky130_fd_sc_hd__buf_1
XFILLER_44_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14592_ _11327_/X _14592_/D VGND VGND VPWR VPWR _14592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13543_ _13542_/X _13086_/X _14337_/Q VGND VGND VPWR VPWR _13543_/X sky130_fd_sc_hd__mux2_1
X_10755_ _10755_/A VGND VGND VPWR VPWR _11506_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13474_ _13473_/X rdata[16] _13516_/S VGND VGND VPWR VPWR _13474_/X sky130_fd_sc_hd__mux2_2
X_10686_ _10783_/A VGND VGND VPWR VPWR _10719_/A sky130_fd_sc_hd__clkbuf_2
X_15213_ _08875_/X _15213_/D VGND VGND VPWR VPWR _15213_/Q sky130_fd_sc_hd__dfxtp_1
X_12425_ _12456_/A _12425_/B VGND VGND VPWR VPWR _12452_/B sky130_fd_sc_hd__or2_1
XFILLER_139_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15144_ _09133_/X _15144_/D VGND VGND VPWR VPWR _15144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12356_ _12363_/A _12395_/B _12355_/Y VGND VGND VPWR VPWR _12431_/B sky130_fd_sc_hd__a21o_1
XFILLER_99_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11307_ _14598_/Q _11303_/X _11191_/X _11304_/X VGND VGND VPWR VPWR _14598_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15075_ _09405_/X _15075_/D VGND VGND VPWR VPWR _15075_/Q sky130_fd_sc_hd__dfxtp_1
X_12287_ _12287_/A _12287_/B VGND VGND VPWR VPWR _12287_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14026_ _14022_/X _14023_/X _14024_/X _14025_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14026_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11238_ _14618_/Q _11232_/X _11104_/X _11233_/X VGND VGND VPWR VPWR _14618_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11169_ _11177_/A VGND VGND VPWR VPWR _11169_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14928_ _10010_/X _14928_/D VGND VGND VPWR VPWR _14928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14859_ _10264_/X _14859_/D VGND VGND VPWR VPWR _14859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07400_ _07402_/A _13535_/X VGND VGND VPWR VPWR _15590_/D sky130_fd_sc_hd__and2_1
X_08380_ _08416_/A VGND VGND VPWR VPWR _08393_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07331_ _07491_/B _07319_/X _07493_/B _07324_/X VGND VGND VPWR VPWR _07333_/B sky130_fd_sc_hd__o22a_1
XFILLER_32_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07262_ _07270_/A VGND VGND VPWR VPWR _07265_/A sky130_fd_sc_hd__clkbuf_2
X_09001_ _09202_/A VGND VGND VPWR VPWR _09068_/A sky130_fd_sc_hd__buf_1
X_07193_ _07254_/B _07177_/B _07188_/X _07190_/Y VGND VGND VPWR VPWR _15663_/D sky130_fd_sc_hd__a211oi_2
XFILLER_145_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09903_ _14953_/Q _09898_/X _09667_/X _09899_/X VGND VGND VPWR VPWR _14953_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09834_ _09836_/A VGND VGND VPWR VPWR _09834_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09765_ _09785_/A VGND VGND VPWR VPWR _09772_/A sky130_fd_sc_hd__buf_1
XFILLER_27_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08716_ _08746_/A VGND VGND VPWR VPWR _08735_/A sky130_fd_sc_hd__buf_1
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09696_ _15011_/Q _09525_/A _09695_/X _09530_/A VGND VGND VPWR VPWR _15011_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08647_ _08647_/A VGND VGND VPWR VPWR _08647_/X sky130_fd_sc_hd__buf_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08578_ _15292_/Q _08576_/X _08390_/X _08577_/X VGND VGND VPWR VPWR _15292_/D sky130_fd_sc_hd__a22o_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07529_ _12019_/A VGND VGND VPWR VPWR _07934_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10540_ _10540_/A VGND VGND VPWR VPWR _10540_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10471_ _14810_/Q _10465_/X _10336_/X _10466_/X VGND VGND VPWR VPWR _14810_/D sky130_fd_sc_hd__a22o_1
X_12210_ _15532_/Q VGND VGND VPWR VPWR _12230_/A sky130_fd_sc_hd__inv_2
X_13190_ _13189_/X _13274_/X _15565_/Q VGND VGND VPWR VPWR _13190_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12141_ _12139_/X _12082_/X _12668_/A _12107_/A VGND VGND VPWR VPWR _12287_/B sky130_fd_sc_hd__o22a_1
XFILLER_150_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12072_ _12128_/A VGND VGND VPWR VPWR _12105_/A sky130_fd_sc_hd__buf_1
XFILLER_150_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11023_ _11023_/A VGND VGND VPWR VPWR _11023_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12974_ _12974_/A _12974_/B _13387_/X VGND VGND VPWR VPWR _13386_/S sky130_fd_sc_hd__or3b_1
XFILLER_92_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14713_ _10873_/X _14713_/D VGND VGND VPWR VPWR _14713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11925_ _11946_/A VGND VGND VPWR VPWR _11925_/X sky130_fd_sc_hd__buf_1
XFILLER_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11856_ _11865_/A VGND VGND VPWR VPWR _11856_/X sky130_fd_sc_hd__buf_1
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14644_ _11129_/X _14644_/D VGND VGND VPWR VPWR _14644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10807_ _10817_/A VGND VGND VPWR VPWR _10807_/X sky130_fd_sc_hd__clkbuf_1
X_14575_ _11388_/X _14575_/D VGND VGND VPWR VPWR _14575_/Q sky130_fd_sc_hd__dfxtp_1
X_11787_ _11807_/A VGND VGND VPWR VPWR _11792_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13526_ _13525_/X _14335_/D _15506_/Q VGND VGND VPWR VPWR _13526_/X sky130_fd_sc_hd__mux2_1
X_10738_ _10738_/A VGND VGND VPWR VPWR _10738_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13457_ _13456_/X _13081_/X _14336_/Q VGND VGND VPWR VPWR _13457_/X sky130_fd_sc_hd__mux2_1
X_10669_ _14754_/Q _10663_/X _10665_/X _10668_/X VGND VGND VPWR VPWR _14754_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12408_ _12415_/A _12407_/A _12412_/A _12407_/Y VGND VGND VPWR VPWR _12409_/A sky130_fd_sc_hd__o22a_2
X_13388_ _12817_/B _12885_/X _13418_/S VGND VGND VPWR VPWR _13388_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12339_ _12699_/B VGND VGND VPWR VPWR _12417_/A sky130_fd_sc_hd__buf_1
X_15127_ _09205_/X _15127_/D VGND VGND VPWR VPWR _15127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15058_ _09470_/X _15058_/D VGND VGND VPWR VPWR _15058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14009_ _14847_/Q _14879_/Q _14911_/Q _14943_/Q _14060_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14009_/X sky130_fd_sc_hd__mux4_2
X_07880_ _07880_/A VGND VGND VPWR VPWR _07880_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_opt_5_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR clkbuf_opt_5_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09550_ _15039_/Q _09544_/X _09546_/X _09549_/X VGND VGND VPWR VPWR _15039_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08501_ _08508_/A VGND VGND VPWR VPWR _08501_/X sky130_fd_sc_hd__clkbuf_1
X_09481_ _15055_/Q _09475_/X _09240_/X _09476_/X VGND VGND VPWR VPWR _15055_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08432_ _14322_/Q VGND VGND VPWR VPWR _10739_/A sky130_fd_sc_hd__buf_1
XFILLER_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08363_ _08374_/A VGND VGND VPWR VPWR _08363_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07314_ _07314_/A _15528_/D VGND VGND VPWR VPWR _15604_/D sky130_fd_sc_hd__nor2b_1
XFILLER_32_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08294_ _08294_/A VGND VGND VPWR VPWR _10270_/A sky130_fd_sc_hd__buf_1
XFILLER_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07245_ _07288_/B _07241_/X _13092_/X _13091_/X _07184_/X VGND VGND VPWR VPWR _15638_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07176_ _07255_/B _07194_/A VGND VGND VPWR VPWR _07177_/B sky130_fd_sc_hd__or2_2
XFILLER_118_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09817_ _09817_/A VGND VGND VPWR VPWR _09822_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09748_ _09768_/A VGND VGND VPWR VPWR _09748_/X sky130_fd_sc_hd__buf_1
XFILLER_74_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09679_ _15015_/Q _09675_/X _09677_/X _09678_/X VGND VGND VPWR VPWR _15015_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11710_ _11712_/A VGND VGND VPWR VPWR _11710_/X sky130_fd_sc_hd__clkbuf_1
X_12690_ _12690_/A _12690_/B VGND VGND VPWR VPWR _12690_/X sky130_fd_sc_hd__and2_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11647_/A VGND VGND VPWR VPWR _11641_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _15669_/CLK pc[21] VGND VGND VPWR VPWR _14360_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _11587_/A VGND VGND VPWR VPWR _11585_/A sky130_fd_sc_hd__buf_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _13369_/X _13365_/X _13408_/S VGND VGND VPWR VPWR _13311_/X sky130_fd_sc_hd__mux2_1
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10523_ _10555_/A VGND VGND VPWR VPWR _10542_/A sky130_fd_sc_hd__buf_2
X_14291_ _14287_/X _14288_/X _14289_/X _14290_/X _14397_/Q _14398_/Q VGND VGND VPWR
+ VPWR _14291_/X sky130_fd_sc_hd__mux4_1
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13242_ _13294_/X _13293_/X _13393_/S VGND VGND VPWR VPWR _13242_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10454_ _10454_/A VGND VGND VPWR VPWR _10516_/A sky130_fd_sc_hd__clkbuf_4
X_13173_ _13177_/X _13187_/X _13415_/S VGND VGND VPWR VPWR _13173_/X sky130_fd_sc_hd__mux2_1
X_10385_ _10492_/A VGND VGND VPWR VPWR _10462_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12124_ _12635_/A _12123_/B _12290_/A VGND VGND VPWR VPWR _12651_/A sky130_fd_sc_hd__a21oi_2
XFILLER_111_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12055_ _12049_/A _12980_/B _12052_/X _12054_/X VGND VGND VPWR VPWR _12055_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_77_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11006_ _11015_/A VGND VGND VPWR VPWR _11006_/X sky130_fd_sc_hd__buf_1
XFILLER_78_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12957_ _12957_/A _12957_/B _12957_/C _12957_/D VGND VGND VPWR VPWR _12959_/A sky130_fd_sc_hd__or4_4
XFILLER_61_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11908_ _11934_/A VGND VGND VPWR VPWR _11919_/A sky130_fd_sc_hd__buf_1
X_12888_ _15530_/Q VGND VGND VPWR VPWR _12888_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_260 _14312_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14627_ _11200_/X _14627_/D VGND VGND VPWR VPWR _14627_/Q sky130_fd_sc_hd__dfxtp_1
X_11839_ _11839_/A VGND VGND VPWR VPWR _11848_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14558_ _11454_/X _14558_/D VGND VGND VPWR VPWR _14558_/Q sky130_fd_sc_hd__dfxtp_1
X_13509_ _13926_/X _13931_/X _13521_/S VGND VGND VPWR VPWR _13509_/X sky130_fd_sc_hd__mux2_2
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14489_ _11721_/X _14489_/D VGND VGND VPWR VPWR _14489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08981_ _15188_/Q _08974_/X _08848_/X _08976_/X VGND VGND VPWR VPWR _15188_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07932_ _07932_/A VGND VGND VPWR VPWR _07932_/X sky130_fd_sc_hd__buf_1
XFILLER_130_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07863_ _07863_/A _07863_/B VGND VGND VPWR VPWR _07864_/C sky130_fd_sc_hd__nand2_1
XFILLER_56_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09602_ _15029_/Q _09593_/X _09601_/X _09597_/X VGND VGND VPWR VPWR _15029_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07794_ _07793_/A _07792_/Y _07793_/Y _07792_/A _07640_/A VGND VGND VPWR VPWR _15458_/D
+ sky130_fd_sc_hd__o221a_1
X_09533_ _10671_/A VGND VGND VPWR VPWR _10303_/A sky130_fd_sc_hd__buf_1
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09464_ _15060_/Q _09456_/X _09220_/X _09458_/X VGND VGND VPWR VPWR _15060_/D sky130_fd_sc_hd__a22o_1
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ _15320_/Q _08405_/X _08414_/X _08409_/X VGND VGND VPWR VPWR _15320_/D sky130_fd_sc_hd__a22o_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09395_ _09395_/A VGND VGND VPWR VPWR _09395_/X sky130_fd_sc_hd__buf_1
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08346_ _10664_/A VGND VGND VPWR VPWR _09153_/A sky130_fd_sc_hd__buf_1
XFILLER_149_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08277_ _08281_/A VGND VGND VPWR VPWR _08277_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07228_ _07228_/A VGND VGND VPWR VPWR _07228_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07159_ _07280_/B _07159_/B VGND VGND VPWR VPWR _07225_/A sky130_fd_sc_hd__or2_1
X_10170_ _14886_/Q _10166_/X _10055_/X _10167_/X VGND VGND VPWR VPWR _14886_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13860_ _14958_/Q _15054_/Q _15022_/Q _15086_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13860_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12811_ _12846_/B _13286_/X VGND VGND VPWR VPWR _12811_/X sky130_fd_sc_hd__or2_1
XFILLER_28_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13791_ _13787_/X _13788_/X _13789_/X _13790_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13791_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15530_ _15578_/CLK _15530_/D VGND VGND VPWR VPWR _15530_/Q sky130_fd_sc_hd__dfxtp_1
X_12742_ _12879_/A _12913_/B _13261_/X _12741_/X VGND VGND VPWR VPWR _12742_/X sky130_fd_sc_hd__o2bb2a_1
X_15461_ _15667_/CLK _15461_/D VGND VGND VPWR VPWR _15461_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _13361_/X _12620_/X _12670_/X _12672_/Y VGND VGND VPWR VPWR _12673_/X sky130_fd_sc_hd__o22a_1
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11643_/A VGND VGND VPWR VPWR _11624_/X sky130_fd_sc_hd__buf_1
X_14412_ _11990_/X _14412_/D VGND VGND VPWR VPWR _14412_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ _08116_/X _15392_/D VGND VGND VPWR VPWR _15392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14343_ _15648_/CLK pc[4] VGND VGND VPWR VPWR _14343_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11555_ _14535_/Q _11552_/X _11553_/X _11554_/X VGND VGND VPWR VPWR _14535_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10506_ _10506_/A VGND VGND VPWR VPWR _10506_/X sky130_fd_sc_hd__buf_1
XFILLER_7_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14274_ _15172_/Q _15140_/Q _14756_/Q _14788_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14274_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11486_ _11493_/A VGND VGND VPWR VPWR _11486_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13225_ _13226_/X _13246_/X _13408_/S VGND VGND VPWR VPWR _13225_/X sky130_fd_sc_hd__mux2_1
X_10437_ _10447_/A VGND VGND VPWR VPWR _10437_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater9 _15563_/Q VGND VGND VPWR VPWR _13408_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13156_ _12570_/X _12570_/A _13157_/S VGND VGND VPWR VPWR _13156_/X sky130_fd_sc_hd__mux2_1
X_10368_ _10380_/A VGND VGND VPWR VPWR _10368_/X sky130_fd_sc_hd__buf_1
X_12107_ _12107_/A VGND VGND VPWR VPWR _12300_/A sky130_fd_sc_hd__buf_1
X_13087_ _12455_/X _15589_/Q _13090_/S VGND VGND VPWR VPWR _13087_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10299_ _10315_/A VGND VGND VPWR VPWR _10300_/A sky130_fd_sc_hd__buf_1
XFILLER_111_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12038_ _15525_/Q _15524_/Q _15528_/Q VGND VGND VPWR VPWR _12039_/C sky130_fd_sc_hd__or3_1
XFILLER_66_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13989_ _14849_/Q _14881_/Q _14913_/Q _14945_/Q _07387_/A _14060_/S1 VGND VGND VPWR
+ VPWR _13989_/X sky130_fd_sc_hd__mux4_2
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15659_ _15663_/CLK _15659_/D VGND VGND VPWR VPWR _15659_/Q sky130_fd_sc_hd__dfxtp_1
X_08200_ _08200_/A VGND VGND VPWR VPWR _08200_/X sky130_fd_sc_hd__clkbuf_1
X_09180_ _09180_/A VGND VGND VPWR VPWR _09180_/X sky130_fd_sc_hd__buf_1
X_08131_ _08161_/A VGND VGND VPWR VPWR _08150_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08062_ _08077_/A VGND VGND VPWR VPWR _08062_/X sky130_fd_sc_hd__buf_1
XFILLER_146_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08964_ _08964_/A VGND VGND VPWR VPWR _08964_/X sky130_fd_sc_hd__buf_1
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07915_ _14301_/Q VGND VGND VPWR VPWR _08925_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_130_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08895_ _09267_/A VGND VGND VPWR VPWR _08895_/X sky130_fd_sc_hd__buf_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07846_ _07846_/A VGND VGND VPWR VPWR _07846_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07777_ _07703_/X _07777_/B _07777_/C _07777_/D VGND VGND VPWR VPWR _07821_/A sky130_fd_sc_hd__and4b_1
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09516_ _15044_/Q _09410_/A _09287_/X _09413_/A VGND VGND VPWR VPWR _15044_/D sky130_fd_sc_hd__a22o_1
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09447_ _15065_/Q _09445_/X _09196_/X _09446_/X VGND VGND VPWR VPWR _15065_/D sky130_fd_sc_hd__a22o_1
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09378_ _15085_/Q _09375_/X _09250_/X _09377_/X VGND VGND VPWR VPWR _15085_/D sky130_fd_sc_hd__a22o_1
XFILLER_12_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08329_ _08357_/A VGND VGND VPWR VPWR _08334_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11340_ _11342_/A VGND VGND VPWR VPWR _11340_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11271_ _11271_/A VGND VGND VPWR VPWR _11278_/A sky130_fd_sc_hd__buf_1
XFILLER_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13010_ _14354_/Q VGND VGND VPWR VPWR _13010_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10222_ _14872_/Q _10217_/X _09977_/X _10218_/X VGND VGND VPWR VPWR _14872_/D sky130_fd_sc_hd__a22o_1
XFILLER_134_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10153_ _10153_/A VGND VGND VPWR VPWR _10153_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14961_ _09874_/X _14961_/D VGND VGND VPWR VPWR _14961_/Q sky130_fd_sc_hd__dfxtp_1
X_10084_ _10084_/A VGND VGND VPWR VPWR _10146_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13912_ _15208_/Q _14536_/Q _14984_/Q _15400_/Q _13945_/S0 _14400_/Q VGND VGND VPWR
+ VPWR _13912_/X sky130_fd_sc_hd__mux4_2
X_14892_ _10151_/X _14892_/D VGND VGND VPWR VPWR _14892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13843_ _14671_/Q _15247_/Q _14735_/Q _14703_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13843_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10986_ _10986_/A VGND VGND VPWR VPWR _10986_/X sky130_fd_sc_hd__buf_1
X_13774_ _15190_/Q _15158_/Q _14774_/Q _14806_/Q _13918_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13774_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15513_ _15527_/CLK _15513_/D VGND VGND VPWR VPWR _15513_/Q sky130_fd_sc_hd__dfxtp_1
X_12725_ _12725_/A VGND VGND VPWR VPWR _12730_/A sky130_fd_sc_hd__buf_2
X_15444_ _15458_/CLK _15444_/D VGND VGND VPWR VPWR data_address[17] sky130_fd_sc_hd__dfxtp_1
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ _12909_/B VGND VGND VPWR VPWR _12656_/Y sky130_fd_sc_hd__inv_2
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ _14523_/Q _11603_/X _11467_/X _11604_/X VGND VGND VPWR VPWR _14523_/D sky130_fd_sc_hd__a22o_1
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15375_ _08176_/X _15375_/D VGND VGND VPWR VPWR _15375_/Q sky130_fd_sc_hd__dfxtp_1
X_12587_ _12586_/A _12586_/B _12585_/Y _12585_/A _12586_/Y VGND VGND VPWR VPWR _12587_/X
+ sky130_fd_sc_hd__o32a_2
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14326_ _14328_/CLK _14326_/D VGND VGND VPWR VPWR _14326_/Q sky130_fd_sc_hd__dfxtp_1
X_11538_ _14539_/Q _11527_/X _11537_/X _11530_/X VGND VGND VPWR VPWR _14539_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14257_ _14630_/Q _14598_/Q _14566_/Q _15366_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14257_/X sky130_fd_sc_hd__mux4_1
X_11469_ _11469_/A VGND VGND VPWR VPWR _11478_/A sky130_fd_sc_hd__buf_1
X_13208_ _13210_/X _13251_/X _13393_/S VGND VGND VPWR VPWR _13208_/X sky130_fd_sc_hd__mux2_1
X_14188_ _14509_/Q _14477_/Q _14445_/Q _14413_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14188_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13139_ _12730_/A _13008_/Y _13152_/S VGND VGND VPWR VPWR _13139_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07700_ _07650_/A _13136_/X _07650_/A _13136_/X VGND VGND VPWR VPWR _07854_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08680_ _08680_/A VGND VGND VPWR VPWR _08743_/A sky130_fd_sc_hd__buf_4
XFILLER_65_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07631_ _07631_/A VGND VGND VPWR VPWR _07634_/A sky130_fd_sc_hd__buf_1
XFILLER_81_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07562_ _07388_/A _15466_/Q _14397_/Q _07539_/Y _07561_/X VGND VGND VPWR VPWR _07562_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_62_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09301_ _09301_/A VGND VGND VPWR VPWR _09301_/X sky130_fd_sc_hd__buf_1
X_07493_ _07495_/A _07493_/B VGND VGND VPWR VPWR _15526_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09232_ _09232_/A VGND VGND VPWR VPWR _09232_/X sky130_fd_sc_hd__buf_1
XFILLER_61_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09163_ _09175_/A VGND VGND VPWR VPWR _09163_/X sky130_fd_sc_hd__buf_1
X_08114_ _08116_/A VGND VGND VPWR VPWR _08114_/X sky130_fd_sc_hd__clkbuf_1
X_09094_ _09094_/A VGND VGND VPWR VPWR _09094_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08045_ _08045_/A VGND VGND VPWR VPWR _08077_/A sky130_fd_sc_hd__buf_1
XFILLER_134_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09996_ _14932_/Q _09985_/X _09995_/X _09988_/X VGND VGND VPWR VPWR _14932_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08947_ _15199_/Q _08943_/X _08799_/X _08946_/X VGND VGND VPWR VPWR _15199_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08878_ _09250_/A VGND VGND VPWR VPWR _08878_/X sky130_fd_sc_hd__buf_1
XFILLER_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07829_ _07838_/A VGND VGND VPWR VPWR _07872_/A sky130_fd_sc_hd__buf_1
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10840_ _10840_/A VGND VGND VPWR VPWR _10840_/X sky130_fd_sc_hd__buf_1
XFILLER_44_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10771_ _11518_/A VGND VGND VPWR VPWR _10771_/X sky130_fd_sc_hd__buf_1
XFILLER_13_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12510_ _12902_/B _12440_/Y _12509_/Y _12466_/Y VGND VGND VPWR VPWR _12510_/X sky130_fd_sc_hd__a31o_1
X_13490_ _13489_/X _13070_/X _14336_/Q VGND VGND VPWR VPWR _13490_/X sky130_fd_sc_hd__mux2_1
X_12441_ _12435_/X _12440_/A _12902_/B _12440_/Y VGND VGND VPWR VPWR _12443_/B sky130_fd_sc_hd__o22a_1
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15160_ _09079_/X _15160_/D VGND VGND VPWR VPWR _15160_/Q sky130_fd_sc_hd__dfxtp_1
X_12372_ _12352_/X _12359_/X _12362_/X _12363_/A VGND VGND VPWR VPWR _12904_/C sky130_fd_sc_hd__o22a_1
XFILLER_125_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14111_ _14107_/X _14108_/X _14109_/X _14110_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14111_/X sky130_fd_sc_hd__mux4_1
X_11323_ _14594_/Q _11319_/X _11065_/X _11322_/X VGND VGND VPWR VPWR _14594_/D sky130_fd_sc_hd__a22o_1
X_15091_ _09355_/X _15091_/D VGND VGND VPWR VPWR _15091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11254_ _11273_/A VGND VGND VPWR VPWR _11254_/X sky130_fd_sc_hd__buf_1
X_14042_ _15227_/Q _14555_/Q _15003_/Q _15419_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14042_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10205_ _14877_/Q _10196_/X _09954_/X _10199_/X VGND VGND VPWR VPWR _14877_/D sky130_fd_sc_hd__a22o_1
X_11185_ _11190_/A VGND VGND VPWR VPWR _11185_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10136_ _10136_/A VGND VGND VPWR VPWR _10136_/X sky130_fd_sc_hd__buf_1
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10067_ _10067_/A VGND VGND VPWR VPWR _10078_/A sky130_fd_sc_hd__buf_1
X_14944_ _09937_/X _14944_/D VGND VGND VPWR VPWR _14944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14875_ _10212_/X _14875_/D VGND VGND VPWR VPWR _14875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13826_ _13822_/X _13823_/X _13824_/X _13825_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13826_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13757_ _14648_/Q _14616_/Q _14584_/Q _15384_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13757_/X sky130_fd_sc_hd__mux4_2
X_10969_ _10999_/A VGND VGND VPWR VPWR _10988_/A sky130_fd_sc_hd__clkbuf_2
X_12708_ _12708_/A VGND VGND VPWR VPWR _12708_/X sky130_fd_sc_hd__buf_1
XFILLER_31_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13688_ _14527_/Q _14495_/Q _14463_/Q _14431_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13688_/X sky130_fd_sc_hd__mux4_2
X_15427_ _15601_/CLK _15427_/D VGND VGND VPWR VPWR data_address[0] sky130_fd_sc_hd__dfxtp_4
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12639_ _12651_/A _12651_/B VGND VGND VPWR VPWR _12641_/B sky130_fd_sc_hd__and2_1
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15358_ _08247_/X _15358_/D VGND VGND VPWR VPWR _15358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14309_ _14311_/CLK _14309_/D VGND VGND VPWR VPWR _14309_/Q sky130_fd_sc_hd__dfxtp_1
X_15289_ _08586_/X _15289_/D VGND VGND VPWR VPWR _15289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09850_ _09854_/A VGND VGND VPWR VPWR _09850_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08801_ _08879_/A VGND VGND VPWR VPWR _08827_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09781_ _09783_/A VGND VGND VPWR VPWR _09781_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08732_ _08732_/A VGND VGND VPWR VPWR _08732_/X sky130_fd_sc_hd__buf_1
XFILLER_38_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08663_ _10838_/B VGND VGND VPWR VPWR _10949_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07614_ _07631_/A VGND VGND VPWR VPWR _07626_/A sky130_fd_sc_hd__buf_1
XFILLER_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08594_ _08605_/A VGND VGND VPWR VPWR _08603_/A sky130_fd_sc_hd__buf_1
XFILLER_54_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07545_ _07545_/A _07545_/B _07545_/C VGND VGND VPWR VPWR _12986_/A sky130_fd_sc_hd__and3_1
X_07476_ _07478_/A _13493_/X VGND VGND VPWR VPWR _15539_/D sky130_fd_sc_hd__and2_1
XFILLER_139_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09215_ _09215_/A VGND VGND VPWR VPWR _09215_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09146_ _09146_/A VGND VGND VPWR VPWR _09158_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09077_ _15161_/Q _09075_/X _08826_/X _09076_/X VGND VGND VPWR VPWR _15161_/D sky130_fd_sc_hd__a22o_1
X_08028_ _08034_/A VGND VGND VPWR VPWR _08028_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09979_ _09993_/A VGND VGND VPWR VPWR _09990_/A sky130_fd_sc_hd__buf_1
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12990_ _07628_/B _13648_/S _07632_/B _07379_/A _12989_/X VGND VGND VPWR VPWR _12990_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11941_ _11941_/A VGND VGND VPWR VPWR _11941_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14660_ _11054_/X _14660_/D VGND VGND VPWR VPWR _14660_/Q sky130_fd_sc_hd__dfxtp_1
X_11872_ _14446_/Q _11865_/X _08042_/A _11866_/X VGND VGND VPWR VPWR _14446_/D sky130_fd_sc_hd__a22o_1
XFILLER_72_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13611_ _13610_/X _13069_/X _14337_/Q VGND VGND VPWR VPWR _13611_/X sky130_fd_sc_hd__mux2_1
X_10823_ _10823_/A VGND VGND VPWR VPWR _11564_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14591_ _11329_/X _14591_/D VGND VGND VPWR VPWR _14591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13542_ _13541_/X _14331_/D _15506_/Q VGND VGND VPWR VPWR _13542_/X sky130_fd_sc_hd__mux2_1
X_10754_ _10754_/A VGND VGND VPWR VPWR _10754_/X sky130_fd_sc_hd__clkbuf_1
X_13473_ _13806_/X _13811_/X _13521_/S VGND VGND VPWR VPWR _13473_/X sky130_fd_sc_hd__mux2_1
X_10685_ _10685_/A VGND VGND VPWR VPWR _10783_/A sky130_fd_sc_hd__buf_4
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15212_ _08882_/X _15212_/D VGND VGND VPWR VPWR _15212_/Q sky130_fd_sc_hd__dfxtp_1
X_12424_ _12874_/A _13395_/X VGND VGND VPWR VPWR _12425_/B sky130_fd_sc_hd__or2_1
XFILLER_138_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15143_ _09135_/X _15143_/D VGND VGND VPWR VPWR _15143_/Q sky130_fd_sc_hd__dfxtp_1
X_12355_ _12355_/A _12395_/B VGND VGND VPWR VPWR _12355_/Y sky130_fd_sc_hd__nor2_4
XFILLER_153_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11306_ _11308_/A VGND VGND VPWR VPWR _11306_/X sky130_fd_sc_hd__clkbuf_1
X_12286_ _12286_/A VGND VGND VPWR VPWR _12286_/Y sky130_fd_sc_hd__inv_2
X_15074_ _09407_/X _15074_/D VGND VGND VPWR VPWR _15074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14025_ _15133_/Q _15357_/Q _15325_/Q _15293_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14025_/X sky130_fd_sc_hd__mux4_2
X_11237_ _11237_/A VGND VGND VPWR VPWR _11237_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11168_ _11168_/A VGND VGND VPWR VPWR _11177_/A sky130_fd_sc_hd__buf_1
X_10119_ _10137_/A VGND VGND VPWR VPWR _10119_/X sky130_fd_sc_hd__buf_1
X_11099_ _11467_/A VGND VGND VPWR VPWR _11099_/X sky130_fd_sc_hd__buf_1
X_14927_ _10015_/X _14927_/D VGND VGND VPWR VPWR _14927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14858_ _10266_/X _14858_/D VGND VGND VPWR VPWR _14858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13809_ _14835_/Q _14867_/Q _14899_/Q _14931_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13809_/X sky130_fd_sc_hd__mux4_2
XFILLER_23_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14789_ _10540_/X _14789_/D VGND VGND VPWR VPWR _14789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07330_ _14392_/Q VGND VGND VPWR VPWR _07493_/B sky130_fd_sc_hd__inv_2
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07261_ _07274_/A VGND VGND VPWR VPWR _07270_/A sky130_fd_sc_hd__clkbuf_2
X_09000_ _09000_/A VGND VGND VPWR VPWR _09202_/A sky130_fd_sc_hd__buf_1
X_07192_ _13118_/X _07190_/Y _07191_/X _07179_/B VGND VGND VPWR VPWR _15664_/D sky130_fd_sc_hd__o211a_1
XFILLER_129_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09902_ _09906_/A VGND VGND VPWR VPWR _09902_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09833_ _14974_/Q _09825_/X _09553_/X _09828_/X VGND VGND VPWR VPWR _14974_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09764_ _09830_/A VGND VGND VPWR VPWR _09785_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08715_ _15254_/Q _08712_/X _08427_/X _08714_/X VGND VGND VPWR VPWR _15254_/D sky130_fd_sc_hd__a22o_1
XFILLER_73_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09695_ _10434_/A VGND VGND VPWR VPWR _09695_/X sky130_fd_sc_hd__buf_1
XFILLER_132_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08646_ _08652_/A VGND VGND VPWR VPWR _08646_/X sky130_fd_sc_hd__clkbuf_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _08588_/A VGND VGND VPWR VPWR _08577_/X sky130_fd_sc_hd__buf_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07528_ _12012_/A VGND VGND VPWR VPWR _12019_/A sky130_fd_sc_hd__buf_1
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07459_ _07459_/A _13463_/X VGND VGND VPWR VPWR _15549_/D sky130_fd_sc_hd__and2_1
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10470_ _10470_/A VGND VGND VPWR VPWR _10470_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09129_ _09161_/A VGND VGND VPWR VPWR _09146_/A sky130_fd_sc_hd__buf_1
XFILLER_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12140_ _15578_/Q VGND VGND VPWR VPWR _12668_/A sky130_fd_sc_hd__inv_2
XFILLER_136_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12071_ _12071_/A VGND VGND VPWR VPWR _12128_/A sky130_fd_sc_hd__inv_2
XFILLER_151_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11022_ _14670_/Q _11015_/X _10776_/X _11016_/X VGND VGND VPWR VPWR _14670_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12973_ _12977_/A _12984_/B _12973_/C VGND VGND VPWR VPWR _12974_/A sky130_fd_sc_hd__and3_1
XFILLER_57_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14712_ _10877_/X _14712_/D VGND VGND VPWR VPWR _14712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11924_ _11985_/A VGND VGND VPWR VPWR _11946_/A sky130_fd_sc_hd__buf_2
XFILLER_82_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14643_ _11132_/X _14643_/D VGND VGND VPWR VPWR _14643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11855_ _11859_/A VGND VGND VPWR VPWR _11855_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10806_ _10821_/A VGND VGND VPWR VPWR _10817_/A sky130_fd_sc_hd__buf_1
X_14574_ _11390_/X _14574_/D VGND VGND VPWR VPWR _14574_/Q sky130_fd_sc_hd__dfxtp_1
X_11786_ _11820_/A VGND VGND VPWR VPWR _11807_/A sky130_fd_sc_hd__buf_1
XFILLER_13_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13525_ _13524_/X _13581_/A1 _13649_/S VGND VGND VPWR VPWR _13525_/X sky130_fd_sc_hd__mux2_1
X_10737_ _14742_/Q _10732_/X _10734_/X _10736_/X VGND VGND VPWR VPWR _14742_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13456_ _13455_/X rdata[22] _13516_/S VGND VGND VPWR VPWR _13456_/X sky130_fd_sc_hd__mux2_2
X_10668_ _10668_/A VGND VGND VPWR VPWR _10668_/X sky130_fd_sc_hd__buf_1
X_12407_ _12407_/A VGND VGND VPWR VPWR _12407_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13387_ _07619_/B _15520_/Q _15519_/Q VGND VGND VPWR VPWR _13387_/X sky130_fd_sc_hd__mux2_1
X_10599_ _10617_/A VGND VGND VPWR VPWR _10599_/X sky130_fd_sc_hd__buf_1
XFILLER_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15126_ _09208_/X _15126_/D VGND VGND VPWR VPWR _15126_/Q sky130_fd_sc_hd__dfxtp_1
X_12338_ _12338_/A _12338_/B VGND VGND VPWR VPWR _12699_/B sky130_fd_sc_hd__or2_2
XFILLER_127_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15057_ _09472_/X _15057_/D VGND VGND VPWR VPWR _15057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12269_ _12264_/X _12802_/A _12267_/X _12268_/X VGND VGND VPWR VPWR _12269_/X sky130_fd_sc_hd__a31o_1
XFILLER_141_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14008_ _14527_/Q _14495_/Q _14463_/Q _14431_/Q _14060_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14008_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08500_ _15307_/Q _08482_/X _08499_/X _08487_/X VGND VGND VPWR VPWR _15307_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09480_ _09484_/A VGND VGND VPWR VPWR _09480_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08431_ _08431_/A VGND VGND VPWR VPWR _08431_/X sky130_fd_sc_hd__clkbuf_1
X_08362_ _15328_/Q _08344_/X _08361_/X _08350_/X VGND VGND VPWR VPWR _15328_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07313_ _07521_/A _07313_/B VGND VGND VPWR VPWR _15528_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08293_ _15344_/Q _08291_/X _08031_/X _08292_/X VGND VGND VPWR VPWR _15344_/D sky130_fd_sc_hd__a22o_1
XFILLER_137_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07244_ _07288_/B _07241_/X _07287_/B _07191_/X _07243_/Y VGND VGND VPWR VPWR _15639_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07175_ _07256_/B _07175_/B VGND VGND VPWR VPWR _07194_/A sky130_fd_sc_hd__or2_1
XFILLER_117_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09816_ _14978_/Q _09812_/X _09527_/X _09815_/X VGND VGND VPWR VPWR _14978_/D sky130_fd_sc_hd__a22o_1
XFILLER_100_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09747_ _09778_/A VGND VGND VPWR VPWR _09768_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09678_ _09678_/A VGND VGND VPWR VPWR _09678_/X sky130_fd_sc_hd__buf_1
XFILLER_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08629_ _08648_/A VGND VGND VPWR VPWR _08629_/X sky130_fd_sc_hd__buf_1
XFILLER_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11649_/A VGND VGND VPWR VPWR _11647_/A sky130_fd_sc_hd__buf_1
XFILLER_52_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ _14531_/Q _11430_/A _11570_/X _11434_/A VGND VGND VPWR VPWR _14531_/D sky130_fd_sc_hd__a22o_1
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13310_ _13311_/X _12459_/B _13393_/S VGND VGND VPWR VPWR _13310_/X sky130_fd_sc_hd__mux2_2
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10522_ _14795_/Q _10515_/X _10403_/X _10517_/X VGND VGND VPWR VPWR _14795_/D sky130_fd_sc_hd__a22o_1
X_14290_ _14947_/Q _15043_/Q _15011_/Q _15075_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14290_/X sky130_fd_sc_hd__mux4_2
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13241_ _12703_/A _12709_/X _15561_/Q VGND VGND VPWR VPWR _13241_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10453_ _10474_/A VGND VGND VPWR VPWR _10453_/X sky130_fd_sc_hd__buf_1
XFILLER_108_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10384_ _14831_/Q _10378_/X _10383_/X _10380_/X VGND VGND VPWR VPWR _14831_/D sky130_fd_sc_hd__a22o_1
X_13172_ _12480_/B _12435_/X _15561_/Q VGND VGND VPWR VPWR _13172_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12123_ _12635_/A _12123_/B VGND VGND VPWR VPWR _12290_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12054_ _07622_/A _12973_/C _12975_/A VGND VGND VPWR VPWR _12054_/X sky130_fd_sc_hd__o21a_1
X_11005_ _11005_/A VGND VGND VPWR VPWR _11005_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12956_ _12518_/B _12955_/B _12955_/Y VGND VGND VPWR VPWR _12957_/B sky130_fd_sc_hd__o21a_1
XFILLER_92_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11907_ _11907_/A VGND VGND VPWR VPWR _11934_/A sky130_fd_sc_hd__buf_2
XFILLER_18_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12887_ _12886_/X _12885_/X _12365_/X _13360_/X _12826_/X VGND VGND VPWR VPWR _12887_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA_250 _12006_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_261 _13516_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14626_ _11204_/X _14626_/D VGND VGND VPWR VPWR _14626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11838_ _14456_/Q _11834_/X _07988_/A _11835_/X VGND VGND VPWR VPWR _14456_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14557_ _11458_/X _14557_/D VGND VGND VPWR VPWR _14557_/Q sky130_fd_sc_hd__dfxtp_1
X_11769_ _11773_/A VGND VGND VPWR VPWR _11769_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_40_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR _15469_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13508_ _13507_/X _13064_/X _14336_/Q VGND VGND VPWR VPWR _13508_/X sky130_fd_sc_hd__mux2_1
X_14488_ _11727_/X _14488_/D VGND VGND VPWR VPWR _14488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13439_ _13438_/X _13087_/X _14336_/Q VGND VGND VPWR VPWR _13439_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15109_ _09283_/X _15109_/D VGND VGND VPWR VPWR _15109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08980_ _08980_/A VGND VGND VPWR VPWR _08980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07931_ _07952_/A VGND VGND VPWR VPWR _07932_/A sky130_fd_sc_hd__buf_1
XFILLER_69_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07862_ _07861_/A _07860_/Y _07861_/Y _07860_/A _07844_/X VGND VGND VPWR VPWR _15442_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09601_ _10359_/A VGND VGND VPWR VPWR _09601_/X sky130_fd_sc_hd__buf_1
XFILLER_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07793_ _07793_/A VGND VGND VPWR VPWR _07793_/Y sky130_fd_sc_hd__inv_2
X_09532_ _09532_/A VGND VGND VPWR VPWR _09532_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09463_ _09465_/A VGND VGND VPWR VPWR _09463_/X sky130_fd_sc_hd__clkbuf_1
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08414_ _09200_/A VGND VGND VPWR VPWR _08414_/X sky130_fd_sc_hd__buf_1
XFILLER_51_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09394_ _09400_/A VGND VGND VPWR VPWR _09394_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08345_ _14335_/Q VGND VGND VPWR VPWR _10664_/A sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_31_clk _14397_/CLK VGND VGND VPWR VPWR _15456_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08276_ _08285_/A VGND VGND VPWR VPWR _08281_/A sky130_fd_sc_hd__buf_1
X_07227_ _07280_/B _07159_/B _07223_/X _07225_/Y VGND VGND VPWR VPWR _15645_/D sky130_fd_sc_hd__a211oi_2
XFILLER_153_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07158_ _07281_/B _07228_/A VGND VGND VPWR VPWR _07159_/B sky130_fd_sc_hd__or2_1
XFILLER_3_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12810_ _12810_/A VGND VGND VPWR VPWR _12821_/A sky130_fd_sc_hd__buf_1
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13790_ _14965_/Q _15061_/Q _15029_/Q _15093_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13790_/X sky130_fd_sc_hd__mux4_2
XFILLER_55_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12741_ _12782_/A VGND VGND VPWR VPWR _12741_/X sky130_fd_sc_hd__buf_1
XFILLER_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15460_ _15604_/CLK _15460_/D VGND VGND VPWR VPWR _15460_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12672_ _12908_/B VGND VGND VPWR VPWR _12672_/Y sky130_fd_sc_hd__inv_2
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _11992_/X _14411_/D VGND VGND VPWR VPWR _14411_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11623_ _11653_/A VGND VGND VPWR VPWR _11643_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _08119_/X _15391_/D VGND VGND VPWR VPWR _15391_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk _14328_/CLK VGND VGND VPWR VPWR _15590_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _15652_/CLK pc[3] VGND VGND VPWR VPWR _14342_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11554_ _11554_/A VGND VGND VPWR VPWR _11554_/X sky130_fd_sc_hd__buf_1
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10505_ _10505_/A VGND VGND VPWR VPWR _10505_/X sky130_fd_sc_hd__buf_1
XFILLER_144_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14273_ _14660_/Q _15236_/Q _14724_/Q _14692_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14273_/X sky130_fd_sc_hd__mux4_2
X_11485_ _14551_/Q _11474_/X _11484_/X _11476_/X VGND VGND VPWR VPWR _14551_/D sky130_fd_sc_hd__a22o_1
X_13224_ _13223_/X _12878_/X _15565_/Q VGND VGND VPWR VPWR _13224_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10436_ _10449_/A VGND VGND VPWR VPWR _10447_/A sky130_fd_sc_hd__buf_1
XFILLER_109_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13155_ _12572_/X _12572_/A _13157_/S VGND VGND VPWR VPWR _13155_/X sky130_fd_sc_hd__mux2_1
X_10367_ _10367_/A VGND VGND VPWR VPWR _10367_/X sky130_fd_sc_hd__buf_1
XFILLER_151_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12106_ _12106_/A VGND VGND VPWR VPWR _12107_/A sky130_fd_sc_hd__buf_1
XFILLER_2_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13086_ _12422_/Y _15588_/Q _13090_/S VGND VGND VPWR VPWR _13086_/X sky130_fd_sc_hd__mux2_1
X_10298_ _10311_/A VGND VGND VPWR VPWR _10315_/A sky130_fd_sc_hd__inv_2
X_12037_ _12037_/A _15526_/Q VGND VGND VPWR VPWR _12037_/X sky130_fd_sc_hd__or2_1
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13988_ _14529_/Q _14497_/Q _14465_/Q _14433_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13988_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12939_ _12736_/A _12737_/B _12914_/C _12724_/X _12730_/B VGND VGND VPWR VPWR _12939_/X
+ sky130_fd_sc_hd__o32a_1
X_15658_ _15662_/CLK _15658_/D VGND VGND VPWR VPWR _15658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14609_ _11269_/X _14609_/D VGND VGND VPWR VPWR _14609_/Q sky130_fd_sc_hd__dfxtp_1
X_15589_ _15589_/CLK _15589_/D VGND VGND VPWR VPWR _15589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_13_clk clkbuf_opt_11_clk/X VGND VGND VPWR VPWR _14395_/CLK sky130_fd_sc_hd__clkbuf_16
X_08130_ _15389_/Q _08122_/X _07963_/X _08125_/X VGND VGND VPWR VPWR _15389_/D sky130_fd_sc_hd__a22o_1
X_08061_ _08067_/A VGND VGND VPWR VPWR _08061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08963_ _08963_/A VGND VGND VPWR VPWR _08963_/X sky130_fd_sc_hd__buf_1
XFILLER_88_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07914_ _14302_/Q VGND VGND VPWR VPWR _11574_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08894_ _08894_/A VGND VGND VPWR VPWR _08894_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07845_ _07705_/A _07843_/Y _07777_/B _07843_/A _07844_/X VGND VGND VPWR VPWR _15446_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07776_ _07849_/A VGND VGND VPWR VPWR _07777_/D sky130_fd_sc_hd__inv_2
X_09515_ _09515_/A VGND VGND VPWR VPWR _09515_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09446_ _09446_/A VGND VGND VPWR VPWR _09446_/X sky130_fd_sc_hd__buf_1
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09377_ _09396_/A VGND VGND VPWR VPWR _09377_/X sky130_fd_sc_hd__buf_1
X_08328_ _08379_/A VGND VGND VPWR VPWR _08357_/A sky130_fd_sc_hd__buf_1
XFILLER_138_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08259_ _15354_/Q _08252_/X _07978_/X _08253_/X VGND VGND VPWR VPWR _15354_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11270_ _14609_/Q _11264_/X _11144_/X _11265_/X VGND VGND VPWR VPWR _14609_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10221_ _10225_/A VGND VGND VPWR VPWR _10221_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10152_ _14892_/Q _10147_/X _10030_/X _10149_/X VGND VGND VPWR VPWR _14892_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14960_ _09876_/X _14960_/D VGND VGND VPWR VPWR _14960_/Q sky130_fd_sc_hd__dfxtp_1
X_10083_ _10093_/A VGND VGND VPWR VPWR _10083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13911_ _13907_/X _13908_/X _13909_/X _13910_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13911_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14891_ _10153_/X _14891_/D VGND VGND VPWR VPWR _14891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13842_ _15215_/Q _14543_/Q _14991_/Q _15407_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13842_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13773_ _14678_/Q _15254_/Q _14742_/Q _14710_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13773_/X sky130_fd_sc_hd__mux4_2
X_10985_ _10985_/A VGND VGND VPWR VPWR _10985_/X sky130_fd_sc_hd__buf_1
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15512_ _15604_/CLK _15512_/D VGND VGND VPWR VPWR _15512_/Q sky130_fd_sc_hd__dfxtp_1
X_12724_ _15542_/Q VGND VGND VPWR VPWR _12724_/X sky130_fd_sc_hd__buf_1
XFILLER_43_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15443_ _15458_/CLK _15443_/D VGND VGND VPWR VPWR data_address[16] sky130_fd_sc_hd__dfxtp_4
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ _12652_/X _12635_/X _12120_/X _12654_/X VGND VGND VPWR VPWR _12909_/B sky130_fd_sc_hd__o22a_1
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11606_ _11608_/A VGND VGND VPWR VPWR _11606_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15374_ _08178_/X _15374_/D VGND VGND VPWR VPWR _15374_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12586_ _12586_/A _12586_/B VGND VGND VPWR VPWR _12586_/Y sky130_fd_sc_hd__nor2_1
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ _14328_/CLK _14325_/D VGND VGND VPWR VPWR _14325_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11537_ _11537_/A VGND VGND VPWR VPWR _11537_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14256_ _14252_/X _14253_/X _14254_/X _14255_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14256_/X sky130_fd_sc_hd__mux4_2
X_11468_ _14555_/Q _11462_/X _11467_/X _11464_/X VGND VGND VPWR VPWR _14555_/D sky130_fd_sc_hd__a22o_1
X_13207_ _12577_/X _12610_/X _13418_/S VGND VGND VPWR VPWR _13207_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10419_ _10419_/A VGND VGND VPWR VPWR _10419_/X sky130_fd_sc_hd__buf_1
X_14187_ _14637_/Q _14605_/Q _14573_/Q _15373_/Q _14268_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14187_/X sky130_fd_sc_hd__mux4_2
X_11399_ _11403_/A VGND VGND VPWR VPWR _11399_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13138_ _12709_/X _13009_/Y _13152_/S VGND VGND VPWR VPWR _13138_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13069_ _12769_/Y _15571_/Q _13076_/S VGND VGND VPWR VPWR _13069_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_clk clkbuf_opt_2_clk/X VGND VGND VPWR VPWR _14393_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07630_ _07630_/A _07630_/B VGND VGND VPWR VPWR _15468_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07561_ _07387_/A _07531_/Y _07366_/A _15469_/Q VGND VGND VPWR VPWR _07561_/X sky130_fd_sc_hd__o22a_1
XFILLER_34_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09300_ _09312_/A VGND VGND VPWR VPWR _09301_/A sky130_fd_sc_hd__buf_1
XFILLER_22_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07492_ _07496_/A VGND VGND VPWR VPWR _07495_/A sky130_fd_sc_hd__buf_1
XFILLER_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09231_ _09239_/A VGND VGND VPWR VPWR _09231_/X sky130_fd_sc_hd__clkbuf_1
X_09162_ _09190_/A VGND VGND VPWR VPWR _09175_/A sky130_fd_sc_hd__buf_1
XFILLER_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08113_ _15394_/Q _08109_/X _07929_/X _08112_/X VGND VGND VPWR VPWR _15394_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09093_ _15156_/Q _09085_/X _08848_/X _09087_/X VGND VGND VPWR VPWR _15156_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08044_ _08052_/A VGND VGND VPWR VPWR _08044_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09995_ _10363_/A VGND VGND VPWR VPWR _09995_/X sky130_fd_sc_hd__buf_1
XFILLER_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08946_ _08964_/A VGND VGND VPWR VPWR _08946_/X sky130_fd_sc_hd__buf_1
XFILLER_131_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08877_ _08904_/A VGND VGND VPWR VPWR _08877_/X sky130_fd_sc_hd__buf_1
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07828_ _07827_/A _07826_/Y _07827_/Y _07826_/A _07810_/X VGND VGND VPWR VPWR _15450_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07759_ _13151_/X _07757_/Y _13151_/X _07757_/Y VGND VGND VPWR VPWR _07760_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10770_ _10770_/A VGND VGND VPWR VPWR _11518_/A sky130_fd_sc_hd__buf_2
X_09429_ _15071_/Q _09425_/X _09170_/X _09428_/X VGND VGND VPWR VPWR _15071_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12440_ _12440_/A VGND VGND VPWR VPWR _12440_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12371_ _12371_/A VGND VGND VPWR VPWR _12371_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14110_ _14965_/Q _15061_/Q _15029_/Q _15093_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14110_/X sky130_fd_sc_hd__mux4_2
X_11322_ _11322_/A VGND VGND VPWR VPWR _11322_/X sky130_fd_sc_hd__buf_1
X_15090_ _09359_/X _15090_/D VGND VGND VPWR VPWR _15090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14041_ _14037_/X _14038_/X _14039_/X _14040_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14041_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11253_ _11283_/A VGND VGND VPWR VPWR _11273_/A sky130_fd_sc_hd__buf_2
XFILLER_141_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10204_ _10206_/A VGND VGND VPWR VPWR _10204_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11184_ _14632_/Q _11173_/X _11183_/X _11175_/X VGND VGND VPWR VPWR _14632_/D sky130_fd_sc_hd__a22o_1
X_10135_ _10141_/A VGND VGND VPWR VPWR _10135_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10066_ _14915_/Q _09927_/A _10065_/X _09931_/A VGND VGND VPWR VPWR _14915_/D sky130_fd_sc_hd__a22o_1
X_14943_ _09940_/X _14943_/D VGND VGND VPWR VPWR _14943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14874_ _10214_/X _14874_/D VGND VGND VPWR VPWR _14874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13825_ _15121_/Q _15345_/Q _15313_/Q _15281_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13825_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13756_ _13752_/X _13753_/X _13754_/X _13755_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13756_/X sky130_fd_sc_hd__mux4_2
X_10968_ _14687_/Q _10964_/X _10684_/X _10967_/X VGND VGND VPWR VPWR _14687_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12707_ _12707_/A VGND VGND VPWR VPWR _12707_/X sky130_fd_sc_hd__buf_2
X_13687_ _14655_/Q _14623_/Q _14591_/Q _15391_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13687_/X sky130_fd_sc_hd__mux4_2
X_10899_ _10899_/A VGND VGND VPWR VPWR _10899_/X sky130_fd_sc_hd__clkbuf_1
X_15426_ _07912_/X _15426_/D VGND VGND VPWR VPWR _15426_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12638_ _12636_/X _12135_/A _12637_/Y _12289_/A VGND VGND VPWR VPWR _12651_/B sky130_fd_sc_hd__a31o_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15357_ _08249_/X _15357_/D VGND VGND VPWR VPWR _15357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ _12569_/A VGND VGND VPWR VPWR _12570_/A sky130_fd_sc_hd__buf_1
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14308_ _15509_/CLK _14308_/D VGND VGND VPWR VPWR _14308_/Q sky130_fd_sc_hd__dfxtp_2
X_15288_ _08590_/X _15288_/D VGND VGND VPWR VPWR _15288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14239_ _14824_/Q _14856_/Q _14888_/Q _14920_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14239_/X sky130_fd_sc_hd__mux4_2
XFILLER_113_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08800_ _08800_/A VGND VGND VPWR VPWR _08879_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09780_ _14989_/Q _09777_/X _09643_/X _09779_/X VGND VGND VPWR VPWR _14989_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08731_ _08731_/A VGND VGND VPWR VPWR _08731_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08662_ _14303_/Q _14302_/Q _08662_/C VGND VGND VPWR VPWR _10838_/B sky130_fd_sc_hd__or3_1
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07613_ _07613_/A VGND VGND VPWR VPWR _07631_/A sky130_fd_sc_hd__buf_1
X_08593_ _15287_/Q _08587_/X _08420_/X _08588_/X VGND VGND VPWR VPWR _15287_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07544_ _07539_/Y _07533_/A _07540_/Y _14402_/Q _07543_/X VGND VGND VPWR VPWR _07545_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_81_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07475_ _07483_/A VGND VGND VPWR VPWR _07478_/A sky130_fd_sc_hd__buf_1
X_09214_ _15126_/Q _09210_/X _09211_/X _09213_/X VGND VGND VPWR VPWR _15126_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09145_ _15140_/Q _09041_/A _08916_/X _09044_/A VGND VGND VPWR VPWR _15140_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09076_ _09076_/A VGND VGND VPWR VPWR _09076_/X sky130_fd_sc_hd__buf_1
X_08027_ _15409_/Q _08014_/X _08026_/X _08017_/X VGND VGND VPWR VPWR _15409_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09978_ _14936_/Q _09972_/X _09977_/X _09974_/X VGND VGND VPWR VPWR _14936_/D sky130_fd_sc_hd__a22o_1
XFILLER_130_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08929_ _08929_/A VGND VGND VPWR VPWR _08929_/X sky130_fd_sc_hd__buf_1
XFILLER_85_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11940_ _14427_/Q _11936_/X _07973_/A _11937_/X VGND VGND VPWR VPWR _14427_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11871_ _11879_/A VGND VGND VPWR VPWR _11871_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13610_ _13609_/X _14314_/D _15506_/Q VGND VGND VPWR VPWR _13610_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10822_ _10830_/A VGND VGND VPWR VPWR _10822_/X sky130_fd_sc_hd__clkbuf_1
X_14590_ _11338_/X _14590_/D VGND VGND VPWR VPWR _14590_/Q sky130_fd_sc_hd__dfxtp_1
X_13541_ _13540_/X _13581_/A1 _13569_/S VGND VGND VPWR VPWR _13541_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10753_ _14739_/Q _10749_/X _10751_/X _10752_/X VGND VGND VPWR VPWR _14739_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13472_ _13471_/X _13076_/X _14336_/Q VGND VGND VPWR VPWR _13472_/X sky130_fd_sc_hd__mux2_1
X_10684_ _11449_/A VGND VGND VPWR VPWR _10684_/X sky130_fd_sc_hd__buf_1
X_15211_ _08886_/X _15211_/D VGND VGND VPWR VPWR _15211_/Q sky130_fd_sc_hd__dfxtp_1
X_12423_ _13408_/S VGND VGND VPWR VPWR _12874_/A sky130_fd_sc_hd__buf_1
XFILLER_138_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15142_ _09140_/X _15142_/D VGND VGND VPWR VPWR _15142_/Q sky130_fd_sc_hd__dfxtp_1
X_12354_ _12352_/X _12298_/X _12362_/A _12301_/A VGND VGND VPWR VPWR _12395_/B sky130_fd_sc_hd__o22a_2
XFILLER_138_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11305_ _14599_/Q _11303_/X _11187_/X _11304_/X VGND VGND VPWR VPWR _14599_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15073_ _09418_/X _15073_/D VGND VGND VPWR VPWR _15073_/Q sky130_fd_sc_hd__dfxtp_1
X_12285_ _12626_/A _12097_/Y _12284_/Y _12109_/Y VGND VGND VPWR VPWR _12286_/A sky130_fd_sc_hd__a31o_1
X_14024_ _15197_/Q _15165_/Q _14781_/Q _14813_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14024_/X sky130_fd_sc_hd__mux4_2
XFILLER_113_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11236_ _14619_/Q _11232_/X _11099_/X _11233_/X VGND VGND VPWR VPWR _14619_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11167_ _14636_/Q _11160_/X _11166_/X _11163_/X VGND VGND VPWR VPWR _14636_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10118_ _10148_/A VGND VGND VPWR VPWR _10137_/A sky130_fd_sc_hd__buf_2
XFILLER_121_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11098_ _11098_/A VGND VGND VPWR VPWR _11098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14926_ _10019_/X _14926_/D VGND VGND VPWR VPWR _14926_/Q sky130_fd_sc_hd__dfxtp_1
X_10049_ _10054_/A VGND VGND VPWR VPWR _10049_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14857_ _10275_/X _14857_/D VGND VGND VPWR VPWR _14857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13808_ _14515_/Q _14483_/Q _14451_/Q _14419_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13808_/X sky130_fd_sc_hd__mux4_2
X_14788_ _10543_/X _14788_/D VGND VGND VPWR VPWR _14788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13739_ _14842_/Q _14874_/Q _14906_/Q _14938_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13739_/X sky130_fd_sc_hd__mux4_2
XFILLER_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07260_ _07260_/A _07260_/B VGND VGND VPWR VPWR _15628_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07191_ _07221_/A VGND VGND VPWR VPWR _07191_/X sky130_fd_sc_hd__buf_1
X_15409_ _08024_/X _15409_/D VGND VGND VPWR VPWR _15409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09901_ _09910_/A VGND VGND VPWR VPWR _09906_/A sky130_fd_sc_hd__buf_1
XFILLER_59_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09832_ _09836_/A VGND VGND VPWR VPWR _09832_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09763_ _09860_/A VGND VGND VPWR VPWR _09830_/A sky130_fd_sc_hd__buf_1
X_08714_ _08733_/A VGND VGND VPWR VPWR _08714_/X sky130_fd_sc_hd__buf_1
XFILLER_39_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09694_ _10831_/A VGND VGND VPWR VPWR _10434_/A sky130_fd_sc_hd__buf_1
XFILLER_67_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08645_ _08671_/A VGND VGND VPWR VPWR _08652_/A sky130_fd_sc_hd__buf_1
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ _08587_/A VGND VGND VPWR VPWR _08576_/X sky130_fd_sc_hd__buf_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07527_ _11973_/A VGND VGND VPWR VPWR _12012_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07458_ _07459_/A _13460_/X VGND VGND VPWR VPWR _15550_/D sky130_fd_sc_hd__and2_1
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07389_ _07512_/B _07322_/X _12568_/A _07373_/X VGND VGND VPWR VPWR _07389_/X sky130_fd_sc_hd__o22a_1
XFILLER_108_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09128_ _15146_/Q _09126_/X _08891_/X _09127_/X VGND VGND VPWR VPWR _15146_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09059_ _09059_/A VGND VGND VPWR VPWR _09064_/A sky130_fd_sc_hd__buf_1
XFILLER_135_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12070_ _15583_/Q VGND VGND VPWR VPWR _12599_/A sky130_fd_sc_hd__inv_2
XFILLER_1_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11021_ _11023_/A VGND VGND VPWR VPWR _11021_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12972_ _12972_/A VGND VGND VPWR VPWR _13421_/S sky130_fd_sc_hd__inv_2
X_14711_ _10879_/X _14711_/D VGND VGND VPWR VPWR _14711_/Q sky130_fd_sc_hd__dfxtp_1
X_11923_ _11923_/A VGND VGND VPWR VPWR _11985_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14642_ _11137_/X _14642_/D VGND VGND VPWR VPWR _14642_/Q sky130_fd_sc_hd__dfxtp_1
X_11854_ _14452_/Q _11844_/X _08011_/A _11846_/X VGND VGND VPWR VPWR _14452_/D sky130_fd_sc_hd__a22o_1
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10805_ _14729_/Q _10797_/X _10804_/X _10800_/X VGND VGND VPWR VPWR _14729_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14573_ _11392_/X _14573_/D VGND VGND VPWR VPWR _14573_/Q sky130_fd_sc_hd__dfxtp_1
X_11785_ _14471_/Q _11783_/X _11553_/X _11784_/X VGND VGND VPWR VPWR _14471_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13524_ _13976_/X _13981_/X _13648_/S VGND VGND VPWR VPWR _13524_/X sky130_fd_sc_hd__mux2_1
X_10736_ _10767_/A VGND VGND VPWR VPWR _10736_/X sky130_fd_sc_hd__buf_1
XFILLER_13_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13455_ _13746_/X _13751_/X _13521_/S VGND VGND VPWR VPWR _13455_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10667_ _10685_/A VGND VGND VPWR VPWR _10668_/A sky130_fd_sc_hd__buf_1
XFILLER_139_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12406_ _15556_/Q VGND VGND VPWR VPWR _12412_/A sky130_fd_sc_hd__buf_1
XFILLER_127_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13386_ _12052_/X _12027_/A _13386_/S VGND VGND VPWR VPWR _13386_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10598_ _10628_/A VGND VGND VPWR VPWR _10617_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15125_ _09215_/X _15125_/D VGND VGND VPWR VPWR _15125_/Q sky130_fd_sc_hd__dfxtp_1
X_12337_ _12337_/A _12337_/B VGND VGND VPWR VPWR _12338_/B sky130_fd_sc_hd__or2_1
XFILLER_5_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15056_ _09474_/X _15056_/D VGND VGND VPWR VPWR _15056_/Q sky130_fd_sc_hd__dfxtp_1
X_12268_ _12805_/A _12239_/B _12239_/X _12247_/Y VGND VGND VPWR VPWR _12268_/X sky130_fd_sc_hd__a22o_1
X_14007_ _14655_/Q _14623_/Q _14591_/Q _15391_/Q _14060_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14007_/X sky130_fd_sc_hd__mux4_2
X_11219_ _11219_/A VGND VGND VPWR VPWR _11283_/A sky130_fd_sc_hd__buf_2
XFILLER_96_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12199_ _12199_/A VGND VGND VPWR VPWR _12199_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14909_ _10093_/X _14909_/D VGND VGND VPWR VPWR _14909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08430_ _15318_/Q _08424_/X _08427_/X _08429_/X VGND VGND VPWR VPWR _15318_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08361_ _09164_/A VGND VGND VPWR VPWR _08361_/X sky130_fd_sc_hd__buf_1
XFILLER_149_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07312_ _07613_/A VGND VGND VPWR VPWR _07521_/A sky130_fd_sc_hd__buf_1
XFILLER_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08292_ _08292_/A VGND VGND VPWR VPWR _08292_/X sky130_fd_sc_hd__buf_1
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07243_ _07240_/A _07241_/X _07287_/B VGND VGND VPWR VPWR _07243_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_149_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07174_ _07258_/B _07197_/A VGND VGND VPWR VPWR _07175_/B sky130_fd_sc_hd__or2_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09815_ _09815_/A VGND VGND VPWR VPWR _09815_/X sky130_fd_sc_hd__buf_1
XFILLER_59_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09746_ _09767_/A VGND VGND VPWR VPWR _09746_/X sky130_fd_sc_hd__buf_1
XFILLER_36_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09677_ _10419_/A VGND VGND VPWR VPWR _09677_/X sky130_fd_sc_hd__buf_1
XFILLER_15_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08628_ _08628_/A VGND VGND VPWR VPWR _08648_/A sky130_fd_sc_hd__buf_1
XFILLER_82_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08559_ _08559_/A VGND VGND VPWR VPWR _08559_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _11570_/A VGND VGND VPWR VPWR _11570_/X sky130_fd_sc_hd__buf_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10521_ _10521_/A VGND VGND VPWR VPWR _10521_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13240_ _13241_/X _13253_/X _15562_/Q VGND VGND VPWR VPWR _13240_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10452_ _10514_/A VGND VGND VPWR VPWR _10474_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13171_ _13170_/X _13250_/X _15565_/Q VGND VGND VPWR VPWR _13171_/X sky130_fd_sc_hd__mux2_1
X_10383_ _10383_/A VGND VGND VPWR VPWR _10383_/X sky130_fd_sc_hd__buf_1
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12122_ _12120_/X _12092_/X _12652_/A _12300_/A VGND VGND VPWR VPWR _12123_/B sky130_fd_sc_hd__o22a_1
XFILLER_117_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12053_ _15519_/Q VGND VGND VPWR VPWR _12973_/C sky130_fd_sc_hd__buf_1
X_11004_ _14676_/Q _10995_/X _10746_/X _10997_/X VGND VGND VPWR VPWR _14676_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12955_ _15561_/Q _12955_/B VGND VGND VPWR VPWR _12955_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11906_ _14435_/Q _11800_/A _08099_/A _11803_/A VGND VGND VPWR VPWR _14435_/D sky130_fd_sc_hd__a22o_1
XFILLER_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12886_ _12926_/A VGND VGND VPWR VPWR _12886_/X sky130_fd_sc_hd__buf_1
XFILLER_93_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_240 _11354_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_251 _12977_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_262 _14375_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14625_ _11212_/X _14625_/D VGND VGND VPWR VPWR _14625_/Q sky130_fd_sc_hd__dfxtp_1
X_11837_ _11837_/A VGND VGND VPWR VPWR _11837_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14556_ _11461_/X _14556_/D VGND VGND VPWR VPWR _14556_/Q sky130_fd_sc_hd__dfxtp_1
X_11768_ _11777_/A VGND VGND VPWR VPWR _11773_/A sky130_fd_sc_hd__buf_1
XFILLER_14_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10719_ _10719_/A VGND VGND VPWR VPWR _10719_/X sky130_fd_sc_hd__buf_1
XFILLER_147_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13507_ _13506_/X rdata[5] _14338_/Q VGND VGND VPWR VPWR _13507_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14487_ _11729_/X _14487_/D VGND VGND VPWR VPWR _14487_/Q sky130_fd_sc_hd__dfxtp_1
X_11699_ _11699_/A VGND VGND VPWR VPWR _11699_/X sky130_fd_sc_hd__clkbuf_1
X_13438_ _13437_/X rdata[28] _13516_/S VGND VGND VPWR VPWR _13438_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13369_ _13371_/X _13370_/X _13415_/S VGND VGND VPWR VPWR _13369_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15108_ _09286_/X _15108_/D VGND VGND VPWR VPWR _15108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07930_ _07947_/A VGND VGND VPWR VPWR _07952_/A sky130_fd_sc_hd__inv_2
X_15039_ _09541_/X _15039_/D VGND VGND VPWR VPWR _15039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07861_ _07861_/A VGND VGND VPWR VPWR _07861_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09600_ _10739_/A VGND VGND VPWR VPWR _10359_/A sky130_fd_sc_hd__buf_1
XFILLER_83_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07792_ _07792_/A VGND VGND VPWR VPWR _07792_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09531_ _15042_/Q _09525_/X _09527_/X _09530_/X VGND VGND VPWR VPWR _15042_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09462_ _15061_/Q _09456_/X _09216_/X _09458_/X VGND VGND VPWR VPWR _15061_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08413_ _10722_/A VGND VGND VPWR VPWR _09200_/A sky130_fd_sc_hd__buf_1
XFILLER_40_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09393_ _09402_/A VGND VGND VPWR VPWR _09400_/A sky130_fd_sc_hd__buf_1
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08344_ _08344_/A VGND VGND VPWR VPWR _08344_/X sky130_fd_sc_hd__buf_1
XFILLER_20_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08275_ _15350_/Q _08272_/X _08000_/X _08274_/X VGND VGND VPWR VPWR _15350_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07226_ _13100_/X _07225_/Y _07221_/X _07161_/B VGND VGND VPWR VPWR _15646_/D sky130_fd_sc_hd__o211a_1
XFILLER_138_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07157_ _07282_/B _07157_/B VGND VGND VPWR VPWR _07228_/A sky130_fd_sc_hd__or2_1
XFILLER_145_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09729_ _09731_/A VGND VGND VPWR VPWR _09729_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12740_ _12740_/A VGND VGND VPWR VPWR _12782_/A sky130_fd_sc_hd__buf_1
XFILLER_55_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12666_/X _12139_/X _12287_/A _12668_/X VGND VGND VPWR VPWR _12908_/B sky130_fd_sc_hd__o22a_1
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14410_ _11995_/X _14410_/D VGND VGND VPWR VPWR _14410_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11642_/A VGND VGND VPWR VPWR _11622_/X sky130_fd_sc_hd__buf_1
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _08127_/X _15390_/D VGND VGND VPWR VPWR _15390_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _15458_/CLK pc[2] VGND VGND VPWR VPWR _14341_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ _11553_/A VGND VGND VPWR VPWR _11553_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10504_ _10510_/A VGND VGND VPWR VPWR _10504_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14272_ _15204_/Q _14532_/Q _14980_/Q _15396_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14272_/X sky130_fd_sc_hd__mux4_2
XFILLER_109_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11484_ _11484_/A VGND VGND VPWR VPWR _11484_/X sky130_fd_sc_hd__buf_1
X_13223_ _13225_/X _13269_/X _13393_/S VGND VGND VPWR VPWR _13223_/X sky130_fd_sc_hd__mux2_1
X_10435_ _14819_/Q _10296_/A _10434_/X _10300_/A VGND VGND VPWR VPWR _14819_/D sky130_fd_sc_hd__a22o_1
XFILLER_124_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13154_ _12573_/X _12573_/A _13157_/S VGND VGND VPWR VPWR _13154_/X sky130_fd_sc_hd__mux2_1
X_10366_ _10378_/A VGND VGND VPWR VPWR _10366_/X sky130_fd_sc_hd__buf_1
XFILLER_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12105_ _12105_/A VGND VGND VPWR VPWR _12106_/A sky130_fd_sc_hd__buf_1
XFILLER_2_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13085_ _12399_/Y _15587_/Q _13090_/S VGND VGND VPWR VPWR _13085_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10297_ _10297_/A VGND VGND VPWR VPWR _10297_/X sky130_fd_sc_hd__buf_1
X_12036_ _12036_/A _12975_/A VGND VGND VPWR VPWR _12982_/A sky130_fd_sc_hd__or2_2
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13987_ _14657_/Q _14625_/Q _14593_/Q _15393_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13987_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12938_ _12752_/X _12758_/B _12958_/A _12934_/X _12937_/X VGND VGND VPWR VPWR _12938_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15657_ _15662_/CLK _15657_/D VGND VGND VPWR VPWR _15657_/Q sky130_fd_sc_hd__dfxtp_1
X_12869_ _12929_/C VGND VGND VPWR VPWR _12869_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14608_ _11272_/X _14608_/D VGND VGND VPWR VPWR _14608_/Q sky130_fd_sc_hd__dfxtp_1
X_15588_ _15589_/CLK _15588_/D VGND VGND VPWR VPWR _15588_/Q sky130_fd_sc_hd__dfxtp_1
X_14539_ _11536_/X _14539_/D VGND VGND VPWR VPWR _14539_/Q sky130_fd_sc_hd__dfxtp_1
X_08060_ _15403_/Q _08046_/X _08059_/X _08050_/X VGND VGND VPWR VPWR _15403_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08962_ _08968_/A VGND VGND VPWR VPWR _08962_/X sky130_fd_sc_hd__clkbuf_1
X_07913_ _14303_/Q VGND VGND VPWR VPWR _08925_/A sky130_fd_sc_hd__clkbuf_1
X_08893_ _15210_/Q _08890_/X _08891_/X _08892_/X VGND VGND VPWR VPWR _15210_/D sky130_fd_sc_hd__a22o_1
X_07844_ _07869_/A VGND VGND VPWR VPWR _07844_/X sky130_fd_sc_hd__buf_1
XFILLER_84_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07775_ _07706_/X _07709_/X _07710_/X _07712_/X _07774_/X VGND VGND VPWR VPWR _07849_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09514_ _15045_/Q _09505_/X _09284_/X _09506_/X VGND VGND VPWR VPWR _15045_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09445_ _09445_/A VGND VGND VPWR VPWR _09445_/X sky130_fd_sc_hd__buf_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09376_ _09376_/A VGND VGND VPWR VPWR _09396_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08327_ _15335_/Q _08325_/X _08079_/X _08326_/X VGND VGND VPWR VPWR _15335_/D sky130_fd_sc_hd__a22o_1
X_08258_ _08260_/A VGND VGND VPWR VPWR _08258_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07209_ _07209_/A VGND VGND VPWR VPWR _07209_/X sky130_fd_sc_hd__buf_1
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08189_ _08189_/A VGND VGND VPWR VPWR _08189_/X sky130_fd_sc_hd__clkbuf_1
X_10220_ _10231_/A VGND VGND VPWR VPWR _10225_/A sky130_fd_sc_hd__buf_2
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10151_ _10153_/A VGND VGND VPWR VPWR _10151_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10082_ _10104_/A VGND VGND VPWR VPWR _10093_/A sky130_fd_sc_hd__buf_1
XFILLER_87_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13910_ _14953_/Q _15049_/Q _15017_/Q _15081_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13910_/X sky130_fd_sc_hd__mux4_1
X_14890_ _10156_/X _14890_/D VGND VGND VPWR VPWR _14890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13841_ _13837_/X _13838_/X _13839_/X _13840_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13841_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13772_ _15222_/Q _14550_/Q _14998_/Q _15414_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13772_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10984_ _10984_/A VGND VGND VPWR VPWR _10984_/X sky130_fd_sc_hd__clkbuf_1
X_15511_ _15604_/CLK _15511_/D VGND VGND VPWR VPWR _15511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12723_ _12684_/X _12722_/X _12684_/X _12722_/X VGND VGND VPWR VPWR _12723_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_31_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15442_ _15458_/CLK _15442_/D VGND VGND VPWR VPWR data_address[15] sky130_fd_sc_hd__dfxtp_1
X_12654_ _15547_/Q VGND VGND VPWR VPWR _12654_/X sky130_fd_sc_hd__buf_1
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11605_ _14524_/Q _11603_/X _11463_/X _11604_/X VGND VGND VPWR VPWR _14524_/D sky130_fd_sc_hd__a22o_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _12585_/A VGND VGND VPWR VPWR _12585_/Y sky130_fd_sc_hd__inv_2
X_15373_ _08181_/X _15373_/D VGND VGND VPWR VPWR _15373_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14324_ _14324_/CLK _14324_/D VGND VGND VPWR VPWR _14324_/Q sky130_fd_sc_hd__dfxtp_1
X_11536_ _11544_/A VGND VGND VPWR VPWR _11536_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14255_ _15110_/Q _15334_/Q _15302_/Q _15270_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14255_/X sky130_fd_sc_hd__mux4_1
X_11467_ _11467_/A VGND VGND VPWR VPWR _11467_/X sky130_fd_sc_hd__buf_1
XFILLER_99_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13206_ _13207_/X _13217_/X _13415_/S VGND VGND VPWR VPWR _13206_/X sky130_fd_sc_hd__mux2_1
X_10418_ _10418_/A VGND VGND VPWR VPWR _10418_/X sky130_fd_sc_hd__buf_1
XFILLER_125_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14186_ _14182_/X _14183_/X _14184_/X _14185_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14186_/X sky130_fd_sc_hd__mux4_2
X_11398_ _11398_/A VGND VGND VPWR VPWR _11403_/A sky130_fd_sc_hd__buf_1
X_13137_ _12703_/A _13010_/Y _13152_/S VGND VGND VPWR VPWR _13137_/X sky130_fd_sc_hd__mux2_1
X_10349_ _10349_/A VGND VGND VPWR VPWR _10349_/X sky130_fd_sc_hd__buf_1
XFILLER_152_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13068_ _12787_/Y _15570_/Q _13076_/S VGND VGND VPWR VPWR _13068_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12019_ _12019_/A VGND VGND VPWR VPWR _12019_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07560_ _07373_/A _07558_/Y _07354_/A _07559_/X VGND VGND VPWR VPWR _07560_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07491_ _07491_/A _07491_/B VGND VGND VPWR VPWR _15527_/D sky130_fd_sc_hd__nor2_1
XFILLER_80_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09230_ _09230_/A VGND VGND VPWR VPWR _09239_/A sky130_fd_sc_hd__buf_1
XFILLER_22_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09161_ _09161_/A VGND VGND VPWR VPWR _09190_/A sky130_fd_sc_hd__clkbuf_2
X_08112_ _08112_/A VGND VGND VPWR VPWR _08112_/X sky130_fd_sc_hd__buf_1
X_09092_ _09094_/A VGND VGND VPWR VPWR _09092_/X sky130_fd_sc_hd__clkbuf_1
X_08043_ _15406_/Q _08029_/X _08042_/X _08032_/X VGND VGND VPWR VPWR _15406_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09994_ _10002_/A VGND VGND VPWR VPWR _09994_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08945_ _09007_/A VGND VGND VPWR VPWR _08964_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08876_ _08876_/A VGND VGND VPWR VPWR _08904_/A sky130_fd_sc_hd__buf_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07827_ _07827_/A VGND VGND VPWR VPWR _07827_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07758_ _15593_/Q VGND VGND VPWR VPWR _07760_/B sky130_fd_sc_hd__inv_2
X_07689_ _07689_/A VGND VGND VPWR VPWR _07689_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09428_ _09446_/A VGND VGND VPWR VPWR _09428_/X sky130_fd_sc_hd__buf_1
X_09359_ _09361_/A VGND VGND VPWR VPWR _09359_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12370_ _12670_/A VGND VGND VPWR VPWR _12371_/A sky130_fd_sc_hd__buf_1
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11321_ _11333_/A VGND VGND VPWR VPWR _11322_/A sky130_fd_sc_hd__buf_1
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14040_ _14972_/Q _15068_/Q _15036_/Q _15100_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _14040_/X sky130_fd_sc_hd__mux4_2
X_11252_ _11260_/A VGND VGND VPWR VPWR _11252_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10203_ _14878_/Q _10196_/X _09950_/X _10199_/X VGND VGND VPWR VPWR _14878_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11183_ _11549_/A VGND VGND VPWR VPWR _11183_/X sky130_fd_sc_hd__buf_1
XFILLER_133_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10134_ _10134_/A VGND VGND VPWR VPWR _10141_/A sky130_fd_sc_hd__buf_1
XFILLER_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10065_ _10434_/A VGND VGND VPWR VPWR _10065_/X sky130_fd_sc_hd__buf_1
X_14942_ _09949_/X _14942_/D VGND VGND VPWR VPWR _14942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14873_ _10216_/X _14873_/D VGND VGND VPWR VPWR _14873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13824_ _15185_/Q _15153_/Q _14769_/Q _14801_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13824_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10967_ _10986_/A VGND VGND VPWR VPWR _10967_/X sky130_fd_sc_hd__buf_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13755_ _15128_/Q _15352_/Q _15320_/Q _15288_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13755_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12706_ _12706_/A VGND VGND VPWR VPWR _12707_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10898_ _14706_/Q _10894_/X _10756_/X _10895_/X VGND VGND VPWR VPWR _14706_/D sky130_fd_sc_hd__a22o_1
X_13686_ _13682_/X _13683_/X _13684_/X _13685_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13686_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15425_ _07934_/X _15425_/D VGND VGND VPWR VPWR _15425_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ _12637_/A VGND VGND VPWR VPWR _12637_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12568_ _12568_/A _12572_/B VGND VGND VPWR VPWR _12568_/Y sky130_fd_sc_hd__nor2_1
X_15356_ _08251_/X _15356_/D VGND VGND VPWR VPWR _15356_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11519_ _14543_/Q _11513_/X _11518_/X _11515_/X VGND VGND VPWR VPWR _14543_/D sky130_fd_sc_hd__a22o_1
X_14307_ _15517_/CLK _14307_/D VGND VGND VPWR VPWR _14307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15287_ _08592_/X _15287_/D VGND VGND VPWR VPWR _15287_/Q sky130_fd_sc_hd__dfxtp_1
X_12499_ _15559_/Q VGND VGND VPWR VPWR _12951_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14238_ _14504_/Q _14472_/Q _14440_/Q _14408_/Q _14238_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14238_/X sky130_fd_sc_hd__mux4_2
XFILLER_113_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14169_ _14831_/Q _14863_/Q _14895_/Q _14927_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14169_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08730_ _15249_/Q _08723_/X _08460_/X _08724_/X VGND VGND VPWR VPWR _15249_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08661_ _11428_/B VGND VGND VPWR VPWR _09408_/A sky130_fd_sc_hd__buf_1
XFILLER_94_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07612_ _07612_/A _13059_/X VGND VGND VPWR VPWR _15474_/D sky130_fd_sc_hd__and2_1
XFILLER_26_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08592_ _08592_/A VGND VGND VPWR VPWR _08592_/X sky130_fd_sc_hd__clkbuf_1
X_07543_ _15467_/Q _07541_/Y _15466_/Q _07542_/Y VGND VGND VPWR VPWR _07543_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07474_ _07573_/A VGND VGND VPWR VPWR _07483_/A sky130_fd_sc_hd__buf_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09213_ _09237_/A VGND VGND VPWR VPWR _09213_/X sky130_fd_sc_hd__buf_1
X_09144_ _09144_/A VGND VGND VPWR VPWR _09144_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09075_ _09075_/A VGND VGND VPWR VPWR _09075_/X sky130_fd_sc_hd__buf_1
XFILLER_135_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08026_ _08026_/A VGND VGND VPWR VPWR _08026_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09977_ _10344_/A VGND VGND VPWR VPWR _09977_/X sky130_fd_sc_hd__buf_1
XFILLER_130_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08928_ _08941_/A VGND VGND VPWR VPWR _08929_/A sky130_fd_sc_hd__buf_1
XFILLER_85_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08859_ _08885_/A VGND VGND VPWR VPWR _08868_/A sky130_fd_sc_hd__buf_1
XFILLER_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11870_ _11870_/A VGND VGND VPWR VPWR _11879_/A sky130_fd_sc_hd__buf_2
XFILLER_44_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10821_ _10821_/A VGND VGND VPWR VPWR _10830_/A sky130_fd_sc_hd__buf_2
XFILLER_26_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10752_ _10767_/A VGND VGND VPWR VPWR _10752_/X sky130_fd_sc_hd__buf_1
X_13540_ _14016_/X _14021_/X _14387_/Q VGND VGND VPWR VPWR _13540_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13471_ _13470_/X rdata[17] _13516_/S VGND VGND VPWR VPWR _13471_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10683_ _10683_/A VGND VGND VPWR VPWR _11449_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12422_ _12349_/X _12411_/X _12413_/Y _12418_/X _12421_/X VGND VGND VPWR VPWR _12422_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_15210_ _08889_/X _15210_/D VGND VGND VPWR VPWR _15210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12353_ _15586_/Q VGND VGND VPWR VPWR _12362_/A sky130_fd_sc_hd__inv_2
X_15141_ _09142_/X _15141_/D VGND VGND VPWR VPWR _15141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11304_ _11304_/A VGND VGND VPWR VPWR _11304_/X sky130_fd_sc_hd__buf_1
X_15072_ _09420_/X _15072_/D VGND VGND VPWR VPWR _15072_/Q sky130_fd_sc_hd__dfxtp_1
X_12284_ _12610_/A _12284_/B VGND VGND VPWR VPWR _12284_/Y sky130_fd_sc_hd__nand2_1
X_14023_ _14685_/Q _15261_/Q _14749_/Q _14717_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14023_/X sky130_fd_sc_hd__mux4_2
XFILLER_107_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11235_ _11237_/A VGND VGND VPWR VPWR _11235_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11166_ _11533_/A VGND VGND VPWR VPWR _11166_/X sky130_fd_sc_hd__buf_1
XFILLER_110_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10117_ _10136_/A VGND VGND VPWR VPWR _10117_/X sky130_fd_sc_hd__buf_1
XFILLER_96_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11097_ _14652_/Q _11094_/X _11095_/X _11096_/X VGND VGND VPWR VPWR _14652_/D sky130_fd_sc_hd__a22o_1
X_14925_ _10022_/X _14925_/D VGND VGND VPWR VPWR _14925_/Q sky130_fd_sc_hd__dfxtp_1
X_10048_ _14920_/Q _10037_/X _10047_/X _10039_/X VGND VGND VPWR VPWR _14920_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14856_ _10277_/X _14856_/D VGND VGND VPWR VPWR _14856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13807_ _14643_/Q _14611_/Q _14579_/Q _15379_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13807_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14787_ _10545_/X _14787_/D VGND VGND VPWR VPWR _14787_/Q sky130_fd_sc_hd__dfxtp_1
X_11999_ _12001_/A VGND VGND VPWR VPWR _11999_/X sky130_fd_sc_hd__clkbuf_1
X_13738_ _14522_/Q _14490_/Q _14458_/Q _14426_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13738_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13669_ _14849_/Q _14881_/Q _14913_/Q _14945_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13669_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15408_ _08028_/X _15408_/D VGND VGND VPWR VPWR _15408_/Q sky130_fd_sc_hd__dfxtp_1
X_07190_ _07190_/A VGND VGND VPWR VPWR _07190_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15339_ _08313_/X _15339_/D VGND VGND VPWR VPWR _15339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09900_ _14954_/Q _09898_/X _09662_/X _09899_/X VGND VGND VPWR VPWR _14954_/D sky130_fd_sc_hd__a22o_1
XFILLER_116_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09831_ _09849_/A VGND VGND VPWR VPWR _09836_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_opt_8_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR clkbuf_opt_8_clk/X sky130_fd_sc_hd__clkbuf_16
X_09762_ _14993_/Q _09756_/X _09622_/X _09757_/X VGND VGND VPWR VPWR _14993_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08713_ _08743_/A VGND VGND VPWR VPWR _08733_/A sky130_fd_sc_hd__clkbuf_2
X_09693_ _09693_/A VGND VGND VPWR VPWR _09693_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08644_ _08644_/A VGND VGND VPWR VPWR _08671_/A sky130_fd_sc_hd__buf_2
XFILLER_66_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08575_ _08581_/A VGND VGND VPWR VPWR _08575_/X sky130_fd_sc_hd__clkbuf_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07526_ _11850_/A VGND VGND VPWR VPWR _11973_/A sky130_fd_sc_hd__buf_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07457_ _07459_/A _13457_/X VGND VGND VPWR VPWR _15551_/D sky130_fd_sc_hd__and2_1
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07388_ _07388_/A VGND VGND VPWR VPWR _12568_/A sky130_fd_sc_hd__buf_1
XFILLER_10_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09127_ _09137_/A VGND VGND VPWR VPWR _09127_/X sky130_fd_sc_hd__buf_1
XFILLER_108_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09058_ _15167_/Q _09054_/X _08799_/X _09057_/X VGND VGND VPWR VPWR _15167_/D sky130_fd_sc_hd__a22o_1
XFILLER_151_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08009_ _08019_/A VGND VGND VPWR VPWR _08009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11020_ _14671_/Q _11015_/X _10771_/X _11016_/X VGND VGND VPWR VPWR _14671_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12971_ _12338_/B _12059_/B _12961_/Y _12970_/X VGND VGND VPWR VPWR _12971_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_73_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14710_ _10882_/X _14710_/D VGND VGND VPWR VPWR _14710_/Q sky130_fd_sc_hd__dfxtp_1
X_11922_ _11932_/A VGND VGND VPWR VPWR _11922_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14641_ _11143_/X _14641_/D VGND VGND VPWR VPWR _14641_/Q sky130_fd_sc_hd__dfxtp_1
X_11853_ _11859_/A VGND VGND VPWR VPWR _11853_/X sky130_fd_sc_hd__buf_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10804_ _11545_/A VGND VGND VPWR VPWR _10804_/X sky130_fd_sc_hd__buf_1
X_11784_ _11784_/A VGND VGND VPWR VPWR _11784_/X sky130_fd_sc_hd__buf_1
X_14572_ _11399_/X _14572_/D VGND VGND VPWR VPWR _14572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13523_ _13522_/X _13059_/X _14336_/Q VGND VGND VPWR VPWR _13523_/X sky130_fd_sc_hd__mux2_1
X_10735_ _10783_/A VGND VGND VPWR VPWR _10767_/A sky130_fd_sc_hd__buf_1
XFILLER_14_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13454_ _13453_/X _13082_/X _14336_/Q VGND VGND VPWR VPWR _13454_/X sky130_fd_sc_hd__mux2_1
X_10666_ _10680_/A VGND VGND VPWR VPWR _10685_/A sky130_fd_sc_hd__inv_2
XFILLER_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12405_ _12403_/X _12298_/X _12414_/A _12301_/A VGND VGND VPWR VPWR _12407_/A sky130_fd_sc_hd__o22a_2
X_13385_ _12211_/X _12838_/X _13418_/S VGND VGND VPWR VPWR _13385_/X sky130_fd_sc_hd__mux2_1
X_10597_ _10616_/A VGND VGND VPWR VPWR _10597_/X sky130_fd_sc_hd__buf_1
XFILLER_5_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15124_ _09219_/X _15124_/D VGND VGND VPWR VPWR _15124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12336_ _12336_/A VGND VGND VPWR VPWR _12336_/X sky130_fd_sc_hd__buf_1
XFILLER_142_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15055_ _09480_/X _15055_/D VGND VGND VPWR VPWR _15055_/Q sky130_fd_sc_hd__dfxtp_1
X_12267_ _12854_/A _12261_/Y _12266_/Y _12254_/Y VGND VGND VPWR VPWR _12267_/X sky130_fd_sc_hd__a31o_1
X_11218_ _11228_/A VGND VGND VPWR VPWR _11218_/X sky130_fd_sc_hd__clkbuf_1
X_14006_ _14002_/X _14003_/X _14004_/X _14005_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14006_/X sky130_fd_sc_hd__mux4_2
X_12198_ _15537_/Q VGND VGND VPWR VPWR _12791_/A sky130_fd_sc_hd__buf_1
XFILLER_68_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11149_ _11149_/A VGND VGND VPWR VPWR _11149_/X sky130_fd_sc_hd__buf_1
XFILLER_96_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14908_ _10096_/X _14908_/D VGND VGND VPWR VPWR _14908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14839_ _10348_/X _14839_/D VGND VGND VPWR VPWR _14839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08360_ _10676_/A VGND VGND VPWR VPWR _09164_/A sky130_fd_sc_hd__buf_1
X_07311_ _15667_/Q VGND VGND VPWR VPWR _07613_/A sky130_fd_sc_hd__buf_1
X_08291_ _08291_/A VGND VGND VPWR VPWR _08291_/X sky130_fd_sc_hd__buf_1
XFILLER_149_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07242_ _07242_/A VGND VGND VPWR VPWR _07287_/B sky130_fd_sc_hd__buf_1
X_07173_ _07259_/B _07173_/B VGND VGND VPWR VPWR _07197_/A sky130_fd_sc_hd__or2_1
XFILLER_9_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09814_ _09826_/A VGND VGND VPWR VPWR _09815_/A sky130_fd_sc_hd__buf_1
XFILLER_100_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09745_ _09776_/A VGND VGND VPWR VPWR _09767_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09676_ _10813_/A VGND VGND VPWR VPWR _10419_/A sky130_fd_sc_hd__buf_1
X_08627_ _08647_/A VGND VGND VPWR VPWR _08627_/X sky130_fd_sc_hd__buf_1
XFILLER_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08558_ _15297_/Q _08552_/X _08355_/X _08555_/X VGND VGND VPWR VPWR _15297_/D sky130_fd_sc_hd__a22o_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07509_ _07510_/A _07509_/B VGND VGND VPWR VPWR _15516_/D sky130_fd_sc_hd__nor2_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08489_ _08489_/A VGND VGND VPWR VPWR _08489_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ _14796_/Q _10515_/X _10399_/X _10517_/X VGND VGND VPWR VPWR _14796_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10451_ _10451_/A VGND VGND VPWR VPWR _10514_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13170_ _13169_/X _13210_/X _13393_/S VGND VGND VPWR VPWR _13170_/X sky130_fd_sc_hd__mux2_1
X_10382_ _10382_/A VGND VGND VPWR VPWR _10382_/X sky130_fd_sc_hd__clkbuf_1
X_12121_ _15579_/Q VGND VGND VPWR VPWR _12652_/A sky130_fd_sc_hd__inv_2
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12052_ _12052_/A VGND VGND VPWR VPWR _12052_/X sky130_fd_sc_hd__buf_1
XFILLER_120_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11003_ _11005_/A VGND VGND VPWR VPWR _11003_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12954_ _15529_/Q VGND VGND VPWR VPWR _12955_/B sky130_fd_sc_hd__buf_1
X_11905_ _11905_/A VGND VGND VPWR VPWR _11905_/X sky130_fd_sc_hd__clkbuf_1
X_12885_ _12885_/A VGND VGND VPWR VPWR _12885_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_230 _09376_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_241 _11526_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_252 _12805_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14624_ _11214_/X _14624_/D VGND VGND VPWR VPWR _14624_/Q sky130_fd_sc_hd__dfxtp_1
X_11836_ _14457_/Q _11834_/X _07983_/A _11835_/X VGND VGND VPWR VPWR _14457_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14555_ _11466_/X _14555_/D VGND VGND VPWR VPWR _14555_/Q sky130_fd_sc_hd__dfxtp_1
X_11767_ _14477_/Q _11764_/X _11528_/X _11766_/X VGND VGND VPWR VPWR _14477_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13506_ _13916_/X _13921_/X _13521_/S VGND VGND VPWR VPWR _13506_/X sky130_fd_sc_hd__mux2_4
X_10718_ _11475_/A VGND VGND VPWR VPWR _10718_/X sky130_fd_sc_hd__buf_1
X_14486_ _11731_/X _14486_/D VGND VGND VPWR VPWR _14486_/Q sky130_fd_sc_hd__dfxtp_1
X_11698_ _14496_/Q _11688_/X _11443_/X _11691_/X VGND VGND VPWR VPWR _14496_/D sky130_fd_sc_hd__a22o_1
X_13437_ _13686_/X _13691_/X _14386_/Q VGND VGND VPWR VPWR _13437_/X sky130_fd_sc_hd__mux2_1
X_10649_ _10649_/A VGND VGND VPWR VPWR _10674_/A sky130_fd_sc_hd__buf_1
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13368_ _13372_/X _13369_/X _13408_/S VGND VGND VPWR VPWR _13368_/X sky130_fd_sc_hd__mux2_1
X_15107_ _09289_/X _15107_/D VGND VGND VPWR VPWR _15107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12319_ _12452_/A VGND VGND VPWR VPWR _12319_/X sky130_fd_sc_hd__buf_1
X_13299_ _13298_/X _13303_/X _13393_/S VGND VGND VPWR VPWR _13299_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15038_ _09551_/X _15038_/D VGND VGND VPWR VPWR _15038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07860_ _07860_/A VGND VGND VPWR VPWR _07860_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07791_ _07660_/X _13121_/X _07660_/X _13121_/X VGND VGND VPWR VPWR _07792_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09530_ _09530_/A VGND VGND VPWR VPWR _09530_/X sky130_fd_sc_hd__buf_1
XFILLER_37_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09461_ _09465_/A VGND VGND VPWR VPWR _09461_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08412_ _14325_/Q VGND VGND VPWR VPWR _10722_/A sky130_fd_sc_hd__buf_1
X_09392_ _15080_/Q _09386_/X _09271_/X _09387_/X VGND VGND VPWR VPWR _15080_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08343_ _08364_/A VGND VGND VPWR VPWR _08344_/A sky130_fd_sc_hd__buf_1
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08274_ _08292_/A VGND VGND VPWR VPWR _08274_/X sky130_fd_sc_hd__buf_1
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07225_ _07225_/A VGND VGND VPWR VPWR _07225_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07156_ _07284_/B _07231_/A VGND VGND VPWR VPWR _07157_/B sky130_fd_sc_hd__or2_2
XFILLER_106_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07989_ _15416_/Q _07981_/X _07988_/X _07984_/X VGND VGND VPWR VPWR _15416_/D sky130_fd_sc_hd__a22o_1
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09728_ _15004_/Q _09726_/X _09564_/X _09727_/X VGND VGND VPWR VPWR _15004_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09659_ _09665_/A VGND VGND VPWR VPWR _09659_/X sky130_fd_sc_hd__clkbuf_1
X_12670_ _12670_/A VGND VGND VPWR VPWR _12670_/X sky130_fd_sc_hd__buf_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11651_/A VGND VGND VPWR VPWR _11642_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14340_ _15669_/CLK pc[1] VGND VGND VPWR VPWR _14340_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ _11552_/A VGND VGND VPWR VPWR _11552_/X sky130_fd_sc_hd__buf_1
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10503_ _10512_/A VGND VGND VPWR VPWR _10510_/A sky130_fd_sc_hd__buf_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11483_ _11493_/A VGND VGND VPWR VPWR _11483_/X sky130_fd_sc_hd__clkbuf_2
X_14271_ _14267_/X _14268_/X _14269_/X _14270_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14271_/X sky130_fd_sc_hd__mux4_1
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13222_ _12634_/X _12635_/X _15561_/Q VGND VGND VPWR VPWR _13222_/X sky130_fd_sc_hd__mux2_1
X_10434_ _10434_/A VGND VGND VPWR VPWR _10434_/X sky130_fd_sc_hd__buf_1
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10365_ _10370_/A VGND VGND VPWR VPWR _10365_/X sky130_fd_sc_hd__clkbuf_1
X_13153_ _12575_/X _12575_/A _13157_/S VGND VGND VPWR VPWR _13153_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12104_ _15582_/Q VGND VGND VPWR VPWR _12618_/A sky130_fd_sc_hd__inv_2
XFILLER_151_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13084_ _12375_/Y _15586_/Q _13090_/S VGND VGND VPWR VPWR _13084_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10296_ _10296_/A VGND VGND VPWR VPWR _10296_/X sky130_fd_sc_hd__buf_1
XFILLER_111_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12035_ _12984_/B _12035_/B VGND VGND VPWR VPWR _12975_/A sky130_fd_sc_hd__or2_2
XFILLER_66_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13986_ _13982_/X _13983_/X _13984_/X _13985_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _13986_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12937_ _12937_/A _12937_/B VGND VGND VPWR VPWR _12937_/X sky130_fd_sc_hd__or2_1
XFILLER_34_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15656_ _15662_/CLK _15656_/D VGND VGND VPWR VPWR _15656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12868_ _12343_/A _12867_/B _12867_/Y VGND VGND VPWR VPWR _12929_/C sky130_fd_sc_hd__a21oi_2
X_14607_ _11276_/X _14607_/D VGND VGND VPWR VPWR _14607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11819_ _14462_/Q _11813_/X _07958_/A _11816_/X VGND VGND VPWR VPWR _14462_/D sky130_fd_sc_hd__a22o_1
X_15587_ _15590_/CLK _15587_/D VGND VGND VPWR VPWR _15587_/Q sky130_fd_sc_hd__dfxtp_1
X_12799_ _12799_/A VGND VGND VPWR VPWR _12839_/B sky130_fd_sc_hd__clkbuf_2
X_14538_ _11539_/X _14538_/D VGND VGND VPWR VPWR _14538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14469_ _11790_/X _14469_/D VGND VGND VPWR VPWR _14469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08961_ _08961_/A VGND VGND VPWR VPWR _08968_/A sky130_fd_sc_hd__buf_1
XFILLER_130_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07912_ _07934_/A VGND VGND VPWR VPWR _07912_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08892_ _08906_/A VGND VGND VPWR VPWR _08892_/X sky130_fd_sc_hd__buf_1
XFILLER_69_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07843_ _07843_/A VGND VGND VPWR VPWR _07843_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07774_ _07863_/A _07861_/A _07774_/C _07856_/A VGND VGND VPWR VPWR _07774_/X sky130_fd_sc_hd__or4_4
XFILLER_83_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09513_ _09515_/A VGND VGND VPWR VPWR _09513_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09444_ _09444_/A VGND VGND VPWR VPWR _09444_/X sky130_fd_sc_hd__clkbuf_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09375_ _09395_/A VGND VGND VPWR VPWR _09375_/X sky130_fd_sc_hd__buf_1
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08326_ _08326_/A VGND VGND VPWR VPWR _08326_/X sky130_fd_sc_hd__buf_1
XFILLER_149_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08257_ _15355_/Q _08252_/X _07973_/X _08253_/X VGND VGND VPWR VPWR _15355_/D sky130_fd_sc_hd__a22o_1
X_07208_ _07208_/A VGND VGND VPWR VPWR _07208_/Y sky130_fd_sc_hd__inv_2
X_08188_ _15372_/Q _08183_/X _08054_/X _08185_/X VGND VGND VPWR VPWR _15372_/D sky130_fd_sc_hd__a22o_1
XFILLER_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07139_ _13105_/X VGND VGND VPWR VPWR _07271_/B sky130_fd_sc_hd__inv_2
XFILLER_106_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10150_ _14893_/Q _10147_/X _10025_/X _10149_/X VGND VGND VPWR VPWR _14893_/D sky130_fd_sc_hd__a22o_1
XFILLER_134_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10081_ _10143_/A VGND VGND VPWR VPWR _10104_/A sky130_fd_sc_hd__buf_2
XFILLER_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13840_ _14960_/Q _15056_/Q _15024_/Q _15088_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13840_/X sky130_fd_sc_hd__mux4_2
XFILLER_63_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13771_ _13767_/X _13768_/X _13769_/X _13770_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13771_/X sky130_fd_sc_hd__mux4_1
X_10983_ _14682_/Q _10976_/X _10713_/X _10977_/X VGND VGND VPWR VPWR _14682_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15510_ _15510_/CLK _15510_/D VGND VGND VPWR VPWR _15510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12722_ _12737_/A _12168_/A _12721_/Y VGND VGND VPWR VPWR _12722_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15441_ _15621_/CLK _15441_/D VGND VGND VPWR VPWR data_address[14] sky130_fd_sc_hd__dfxtp_4
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ _12652_/X _12635_/X _12336_/A _13344_/X _12319_/X VGND VGND VPWR VPWR _12653_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ _11613_/A VGND VGND VPWR VPWR _11604_/X sky130_fd_sc_hd__buf_1
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ _08187_/X _15372_/D VGND VGND VPWR VPWR _15372_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _12598_/A _12598_/B VGND VGND VPWR VPWR _12586_/B sky130_fd_sc_hd__and2_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ _15469_/CLK _14323_/D VGND VGND VPWR VPWR _14323_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11535_ _11547_/A VGND VGND VPWR VPWR _11544_/A sky130_fd_sc_hd__buf_1
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14254_ _15174_/Q _15142_/Q _14758_/Q _14790_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14254_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11466_ _11466_/A VGND VGND VPWR VPWR _11466_/X sky130_fd_sc_hd__clkbuf_1
X_13205_ _13206_/X _13226_/X _13408_/S VGND VGND VPWR VPWR _13205_/X sky130_fd_sc_hd__mux2_1
X_10417_ _10422_/A VGND VGND VPWR VPWR _10417_/X sky130_fd_sc_hd__clkbuf_1
X_11397_ _14573_/Q _11394_/X _11161_/X _11396_/X VGND VGND VPWR VPWR _14573_/D sky130_fd_sc_hd__a22o_1
X_14185_ _15117_/Q _15341_/Q _15309_/Q _15277_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14185_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13136_ _12662_/X _13011_/Y _13152_/S VGND VGND VPWR VPWR _13136_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10348_ _10358_/A VGND VGND VPWR VPWR _10348_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13067_ _12795_/Y _15569_/Q _13076_/S VGND VGND VPWR VPWR _13067_/X sky130_fd_sc_hd__mux2_2
X_10279_ _10279_/A VGND VGND VPWR VPWR _10279_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12018_ _12019_/A VGND VGND VPWR VPWR _12018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13969_ _14819_/Q _14851_/Q _14883_/Q _14915_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13969_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07490_ _07517_/A _13523_/X VGND VGND VPWR VPWR _15529_/D sky130_fd_sc_hd__and2_1
XFILLER_34_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15639_ _15669_/CLK _15639_/D VGND VGND VPWR VPWR _15639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09160_ _15137_/Q _09152_/X _09159_/X _09156_/X VGND VGND VPWR VPWR _15137_/D sky130_fd_sc_hd__a22o_1
X_08111_ _08123_/A VGND VGND VPWR VPWR _08112_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09091_ _15157_/Q _09085_/X _08844_/X _09087_/X VGND VGND VPWR VPWR _15157_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_08042_ _08042_/A VGND VGND VPWR VPWR _08042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09993_ _09993_/A VGND VGND VPWR VPWR _10002_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08944_ _08944_/A VGND VGND VPWR VPWR _09007_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08875_ _08882_/A VGND VGND VPWR VPWR _08875_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07826_ _07826_/A VGND VGND VPWR VPWR _07826_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07757_ _15594_/Q VGND VGND VPWR VPWR _07757_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07688_ _13130_/X VGND VGND VPWR VPWR _07688_/X sky130_fd_sc_hd__buf_1
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09427_ _09487_/A VGND VGND VPWR VPWR _09446_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09358_ _15091_/Q _09356_/X _09224_/X _09357_/X VGND VGND VPWR VPWR _15091_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08309_ _15341_/Q _08306_/X _08048_/X _08308_/X VGND VGND VPWR VPWR _15341_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09289_ _09289_/A VGND VGND VPWR VPWR _09289_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11320_ _11330_/A VGND VGND VPWR VPWR _11333_/A sky130_fd_sc_hd__inv_2
XFILLER_126_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11251_ _11271_/A VGND VGND VPWR VPWR _11260_/A sky130_fd_sc_hd__buf_1
XFILLER_153_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10202_ _10206_/A VGND VGND VPWR VPWR _10202_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11182_ _11190_/A VGND VGND VPWR VPWR _11182_/X sky130_fd_sc_hd__clkbuf_1
X_10133_ _14897_/Q _10127_/X _10008_/X _10128_/X VGND VGND VPWR VPWR _14897_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10064_ _10064_/A VGND VGND VPWR VPWR _10064_/X sky130_fd_sc_hd__clkbuf_1
X_14941_ _09953_/X _14941_/D VGND VGND VPWR VPWR _14941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14872_ _10221_/X _14872_/D VGND VGND VPWR VPWR _14872_/Q sky130_fd_sc_hd__dfxtp_1
X_13823_ _14673_/Q _15249_/Q _14737_/Q _14705_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13823_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13754_ _15192_/Q _15160_/Q _14776_/Q _14808_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13754_/X sky130_fd_sc_hd__mux4_2
X_10966_ _11026_/A VGND VGND VPWR VPWR _10986_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12705_ _12460_/X _12691_/Y _12696_/Y _12704_/X VGND VGND VPWR VPWR _12705_/Y sky130_fd_sc_hd__o211ai_2
X_13685_ _15135_/Q _15359_/Q _15327_/Q _15295_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13685_/X sky130_fd_sc_hd__mux4_1
X_10897_ _10899_/A VGND VGND VPWR VPWR _10897_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15424_ _07942_/X _15424_/D VGND VGND VPWR VPWR _15424_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ _12636_/A VGND VGND VPWR VPWR _12636_/X sky130_fd_sc_hd__buf_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ _08256_/X _15355_/D VGND VGND VPWR VPWR _15355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12567_ _12575_/B VGND VGND VPWR VPWR _12572_/B sky130_fd_sc_hd__buf_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14306_ _15469_/CLK _14306_/D VGND VGND VPWR VPWR _14306_/Q sky130_fd_sc_hd__dfxtp_1
X_11518_ _11518_/A VGND VGND VPWR VPWR _11518_/X sky130_fd_sc_hd__buf_1
X_15286_ _08595_/X _15286_/D VGND VGND VPWR VPWR _15286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12498_ _15591_/Q VGND VGND VPWR VPWR _12498_/X sky130_fd_sc_hd__clkbuf_2
X_14237_ _14632_/Q _14600_/Q _14568_/Q _15368_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14237_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11449_ _11449_/A VGND VGND VPWR VPWR _11449_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14168_ _14511_/Q _14479_/Q _14447_/Q _14415_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14168_/X sky130_fd_sc_hd__mux4_2
XFILLER_3_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13119_ _15665_/Q data_address[30] _15667_/Q VGND VGND VPWR VPWR _13119_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14099_ _14838_/Q _14870_/Q _14902_/Q _14934_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14099_/X sky130_fd_sc_hd__mux4_2
XFILLER_100_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08660_ _08660_/A VGND VGND VPWR VPWR _11428_/B sky130_fd_sc_hd__buf_1
XFILLER_94_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07611_ _07638_/A _13060_/X VGND VGND VPWR VPWR _15475_/D sky130_fd_sc_hd__and2_1
X_08591_ _15288_/Q _08587_/X _08414_/X _08588_/X VGND VGND VPWR VPWR _15288_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07542_ _07542_/A VGND VGND VPWR VPWR _07542_/Y sky130_fd_sc_hd__inv_2
X_07473_ _07473_/A VGND VGND VPWR VPWR _07573_/A sky130_fd_sc_hd__buf_1
XFILLER_61_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09212_ _09251_/A VGND VGND VPWR VPWR _09237_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09143_ _15141_/Q _09136_/X _08913_/X _09137_/X VGND VGND VPWR VPWR _15141_/D sky130_fd_sc_hd__a22o_1
X_09074_ _09074_/A VGND VGND VPWR VPWR _09074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08025_ _14318_/Q VGND VGND VPWR VPWR _08026_/A sky130_fd_sc_hd__buf_1
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09976_ _09976_/A VGND VGND VPWR VPWR _09976_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08927_ _10294_/A _10438_/B VGND VGND VPWR VPWR _08941_/A sky130_fd_sc_hd__or2_2
XFILLER_131_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08858_ _08858_/A VGND VGND VPWR VPWR _08885_/A sky130_fd_sc_hd__buf_2
X_07809_ _07809_/A VGND VGND VPWR VPWR _07869_/A sky130_fd_sc_hd__buf_1
XFILLER_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08789_ _09159_/A VGND VGND VPWR VPWR _08789_/X sky130_fd_sc_hd__buf_1
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10820_ _14726_/Q _10812_/X _10819_/X _10815_/X VGND VGND VPWR VPWR _14726_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10751_ _11502_/A VGND VGND VPWR VPWR _10751_/X sky130_fd_sc_hd__buf_1
XFILLER_25_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13470_ _13796_/X _13801_/X _13521_/S VGND VGND VPWR VPWR _13470_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10682_ _10716_/A VGND VGND VPWR VPWR _10682_/X sky130_fd_sc_hd__buf_1
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12421_ _12368_/X _12400_/X _12371_/X _12420_/Y VGND VGND VPWR VPWR _12421_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15140_ _09144_/X _15140_/D VGND VGND VPWR VPWR _15140_/Q sky130_fd_sc_hd__dfxtp_1
X_12352_ _15586_/Q VGND VGND VPWR VPWR _12352_/X sky130_fd_sc_hd__buf_1
X_11303_ _11303_/A VGND VGND VPWR VPWR _11303_/X sky130_fd_sc_hd__buf_1
X_15071_ _09422_/X _15071_/D VGND VGND VPWR VPWR _15071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12283_ _12177_/Y _12209_/X _12747_/A _12282_/X VGND VGND VPWR VPWR _12637_/A sky130_fd_sc_hd__o31a_2
X_14022_ _15229_/Q _14557_/Q _15005_/Q _15421_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14022_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11234_ _14620_/Q _11232_/X _11095_/X _11233_/X VGND VGND VPWR VPWR _14620_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11165_ _11165_/A VGND VGND VPWR VPWR _11165_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10116_ _10146_/A VGND VGND VPWR VPWR _10136_/A sky130_fd_sc_hd__buf_2
X_11096_ _11109_/A VGND VGND VPWR VPWR _11096_/X sky130_fd_sc_hd__buf_1
XFILLER_122_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14924_ _10029_/X _14924_/D VGND VGND VPWR VPWR _14924_/Q sky130_fd_sc_hd__dfxtp_1
X_10047_ _10415_/A VGND VGND VPWR VPWR _10047_/X sky130_fd_sc_hd__buf_1
XFILLER_75_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14855_ _10279_/X _14855_/D VGND VGND VPWR VPWR _14855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13806_ _13802_/X _13803_/X _13804_/X _13805_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13806_/X sky130_fd_sc_hd__mux4_2
X_14786_ _10547_/X _14786_/D VGND VGND VPWR VPWR _14786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11998_ _14410_/Q _11996_/X _08064_/A _11997_/X VGND VGND VPWR VPWR _14410_/D sky130_fd_sc_hd__a22o_1
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13737_ _14650_/Q _14618_/Q _14586_/Q _15386_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13737_/X sky130_fd_sc_hd__mux4_2
X_10949_ _10949_/A _11062_/B VGND VGND VPWR VPWR _10962_/A sky130_fd_sc_hd__or2_2
XFILLER_149_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13668_ _14529_/Q _14497_/Q _14465_/Q _14433_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13668_/X sky130_fd_sc_hd__mux4_1
X_15407_ _08034_/X _15407_/D VGND VGND VPWR VPWR _15407_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12619_ _12610_/X _12618_/X _12416_/X _13209_/X _12417_/X VGND VGND VPWR VPWR _12619_/X
+ sky130_fd_sc_hd__o32a_2
X_13599_ _13598_/X _13072_/X _14337_/Q VGND VGND VPWR VPWR _13599_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15338_ _08315_/X _15338_/D VGND VGND VPWR VPWR _15338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_0 data_address[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15269_ _08652_/X _15269_/D VGND VGND VPWR VPWR _15269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09830_ _09830_/A VGND VGND VPWR VPWR _09849_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09761_ _09761_/A VGND VGND VPWR VPWR _09761_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08712_ _08732_/A VGND VGND VPWR VPWR _08712_/X sky130_fd_sc_hd__buf_1
XFILLER_67_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09692_ _15012_/Q _09525_/A _09691_/X _09530_/A VGND VGND VPWR VPWR _15012_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08643_ _15272_/Q _08637_/X _08517_/X _08638_/X VGND VGND VPWR VPWR _15272_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08574_ _08574_/A VGND VGND VPWR VPWR _08581_/A sky130_fd_sc_hd__buf_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07525_ _11559_/A VGND VGND VPWR VPWR _11850_/A sky130_fd_sc_hd__buf_1
XFILLER_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07456_ _07456_/A VGND VGND VPWR VPWR _07459_/A sky130_fd_sc_hd__clkbuf_1
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07387_ _07387_/A VGND VGND VPWR VPWR _07388_/A sky130_fd_sc_hd__inv_2
XFILLER_148_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09126_ _09136_/A VGND VGND VPWR VPWR _09126_/X sky130_fd_sc_hd__buf_1
XFILLER_108_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09057_ _09076_/A VGND VGND VPWR VPWR _09057_/X sky130_fd_sc_hd__buf_1
XFILLER_135_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08008_ _08023_/A VGND VGND VPWR VPWR _08019_/A sky130_fd_sc_hd__buf_1
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09959_ _09974_/A VGND VGND VPWR VPWR _09959_/X sky130_fd_sc_hd__buf_1
XFILLER_103_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12970_ _12325_/B _12338_/B _12972_/A _12966_/Y _12969_/X VGND VGND VPWR VPWR _12970_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11921_ _11934_/A VGND VGND VPWR VPWR _11932_/A sky130_fd_sc_hd__buf_1
XFILLER_73_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14640_ _11146_/X _14640_/D VGND VGND VPWR VPWR _14640_/Q sky130_fd_sc_hd__dfxtp_1
X_11852_ _11870_/A VGND VGND VPWR VPWR _11859_/A sky130_fd_sc_hd__buf_1
XFILLER_14_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10803_ _10803_/A VGND VGND VPWR VPWR _11545_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14571_ _11401_/X _14571_/D VGND VGND VPWR VPWR _14571_/Q sky130_fd_sc_hd__dfxtp_1
X_11783_ _11783_/A VGND VGND VPWR VPWR _11783_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_52_clk _14315_/CLK VGND VGND VPWR VPWR _15668_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13522_ _13521_/X rdata[0] _14338_/Q VGND VGND VPWR VPWR _13522_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10734_ _11489_/A VGND VGND VPWR VPWR _10734_/X sky130_fd_sc_hd__buf_1
XFILLER_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13453_ _13452_/X rdata[23] _13516_/S VGND VGND VPWR VPWR _13453_/X sky130_fd_sc_hd__mux2_1
X_10665_ _11431_/A VGND VGND VPWR VPWR _10665_/X sky130_fd_sc_hd__clkbuf_2
X_12404_ _15588_/Q VGND VGND VPWR VPWR _12414_/A sky130_fd_sc_hd__inv_2
X_13384_ _12847_/A _12820_/X _13418_/S VGND VGND VPWR VPWR _13384_/X sky130_fd_sc_hd__mux2_1
X_10596_ _10626_/A VGND VGND VPWR VPWR _10616_/A sky130_fd_sc_hd__clkbuf_2
X_15123_ _09222_/X _15123_/D VGND VGND VPWR VPWR _15123_/Q sky130_fd_sc_hd__dfxtp_1
X_12335_ _12739_/A VGND VGND VPWR VPWR _12336_/A sky130_fd_sc_hd__buf_1
XFILLER_5_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15054_ _09482_/X _15054_/D VGND VGND VPWR VPWR _15054_/Q sky130_fd_sc_hd__dfxtp_1
X_12266_ _12836_/A _12266_/B VGND VGND VPWR VPWR _12266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14005_ _15135_/Q _15359_/Q _15327_/Q _15295_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14005_/X sky130_fd_sc_hd__mux4_1
X_11217_ _11239_/A VGND VGND VPWR VPWR _11228_/A sky130_fd_sc_hd__buf_1
XFILLER_96_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12197_ _12195_/X _12081_/A _12788_/A _12130_/A VGND VGND VPWR VPWR _12199_/A sky130_fd_sc_hd__o22a_1
XFILLER_96_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11148_ _11514_/A VGND VGND VPWR VPWR _11148_/X sky130_fd_sc_hd__buf_1
XFILLER_1_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11079_ _11159_/A VGND VGND VPWR VPWR _11107_/A sky130_fd_sc_hd__buf_2
XFILLER_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14907_ _10100_/X _14907_/D VGND VGND VPWR VPWR _14907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14838_ _10351_/X _14838_/D VGND VGND VPWR VPWR _14838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14769_ _10613_/X _14769_/D VGND VGND VPWR VPWR _14769_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_43_clk clkbuf_opt_8_clk/X VGND VGND VPWR VPWR _15597_/CLK sky130_fd_sc_hd__clkbuf_16
X_07310_ _07313_/B _07314_/A VGND VGND VPWR VPWR _07310_/Y sky130_fd_sc_hd__nor2_8
X_08290_ _08290_/A VGND VGND VPWR VPWR _08290_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07241_ _07246_/B VGND VGND VPWR VPWR _07241_/X sky130_fd_sc_hd__buf_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07172_ _07260_/B _07202_/A VGND VGND VPWR VPWR _07173_/B sky130_fd_sc_hd__or2_2
XFILLER_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09813_ _09823_/A VGND VGND VPWR VPWR _09826_/A sky130_fd_sc_hd__inv_2
XFILLER_141_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09744_ _09752_/A VGND VGND VPWR VPWR _09744_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09675_ _09675_/A VGND VGND VPWR VPWR _09675_/X sky130_fd_sc_hd__buf_1
XFILLER_55_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08626_ _08626_/A VGND VGND VPWR VPWR _08647_/A sky130_fd_sc_hd__buf_1
XFILLER_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _08559_/A VGND VGND VPWR VPWR _08557_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_clk _14315_/CLK VGND VGND VPWR VPWR _15510_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07508_ _07510_/A _07508_/B VGND VGND VPWR VPWR _15517_/D sky130_fd_sc_hd__nor2_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08488_ _15309_/Q _08482_/X _08485_/X _08487_/X VGND VGND VPWR VPWR _15309_/D sky130_fd_sc_hd__a22o_1
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07439_ _07443_/A VGND VGND VPWR VPWR _07442_/A sky130_fd_sc_hd__clkbuf_1
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10450_ _10460_/A VGND VGND VPWR VPWR _10450_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09109_ _09120_/A VGND VGND VPWR VPWR _09114_/A sky130_fd_sc_hd__buf_1
X_10381_ _14832_/Q _10378_/X _10379_/X _10380_/X VGND VGND VPWR VPWR _14832_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12120_ _15579_/Q VGND VGND VPWR VPWR _12120_/X sky130_fd_sc_hd__buf_1
XFILLER_151_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12051_ _15526_/Q _12983_/C _15527_/Q VGND VGND VPWR VPWR _12052_/A sky130_fd_sc_hd__or3b_2
XFILLER_117_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11002_ _14677_/Q _10995_/X _10740_/X _10997_/X VGND VGND VPWR VPWR _14677_/D sky130_fd_sc_hd__a22o_1
XFILLER_77_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12953_ _12519_/A _12888_/X _12886_/X _12885_/A VGND VGND VPWR VPWR _12957_/A sky130_fd_sc_hd__o22a_1
XFILLER_46_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11904_ _14436_/Q _11800_/A _08095_/A _11803_/A VGND VGND VPWR VPWR _14436_/D sky130_fd_sc_hd__a22o_1
X_15672_ _15672_/D _12993_/Y VGND VGND VPWR VPWR _15672_/Q sky130_fd_sc_hd__dlxtn_1
X_12884_ _12884_/A VGND VGND VPWR VPWR _12884_/X sky130_fd_sc_hd__buf_1
XANTENNA_220 _15451_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_231 _09487_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_242 _11587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14623_ _11218_/X _14623_/D VGND VGND VPWR VPWR _14623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_253 _12825_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11835_ _11835_/A VGND VGND VPWR VPWR _11835_/X sky130_fd_sc_hd__buf_1
XFILLER_26_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14554_ _11470_/X _14554_/D VGND VGND VPWR VPWR _14554_/Q sky130_fd_sc_hd__dfxtp_1
X_11766_ _11784_/A VGND VGND VPWR VPWR _11766_/X sky130_fd_sc_hd__buf_1
X_13505_ _13504_/X _13065_/X _14336_/Q VGND VGND VPWR VPWR _13505_/X sky130_fd_sc_hd__mux2_1
X_10717_ _10717_/A VGND VGND VPWR VPWR _11475_/A sky130_fd_sc_hd__buf_1
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14485_ _11738_/X _14485_/D VGND VGND VPWR VPWR _14485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11697_ _11699_/A VGND VGND VPWR VPWR _11697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13436_ _13435_/X _13088_/X _14336_/Q VGND VGND VPWR VPWR _13436_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10648_ _14759_/Q _10646_/X _10419_/X _10647_/X VGND VGND VPWR VPWR _14759_/D sky130_fd_sc_hd__a22o_1
XFILLER_127_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13367_ _12395_/A _12388_/X _13418_/S VGND VGND VPWR VPWR _13367_/X sky130_fd_sc_hd__mux2_1
X_10579_ _10583_/A VGND VGND VPWR VPWR _10579_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15106_ _09293_/X _15106_/D VGND VGND VPWR VPWR _15106_/Q sky130_fd_sc_hd__dfxtp_1
X_12318_ _12367_/A VGND VGND VPWR VPWR _12452_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_114_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13298_ _13353_/X _13352_/X _13408_/S VGND VGND VPWR VPWR _13298_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15037_ _09557_/X _15037_/D VGND VGND VPWR VPWR _15037_/Q sky130_fd_sc_hd__dfxtp_1
X_12249_ _15534_/Q VGND VGND VPWR VPWR _12254_/A sky130_fd_sc_hd__inv_2
XFILLER_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07790_ _07659_/X _13122_/X _07789_/Y VGND VGND VPWR VPWR _07793_/A sky130_fd_sc_hd__o21ai_1
XFILLER_68_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09460_ _09469_/A VGND VGND VPWR VPWR _09465_/A sky130_fd_sc_hd__buf_1
XFILLER_52_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08411_ _08411_/A VGND VGND VPWR VPWR _08411_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09391_ _09391_/A VGND VGND VPWR VPWR _09391_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_16_clk _14328_/CLK VGND VGND VPWR VPWR _15498_/CLK sky130_fd_sc_hd__clkbuf_16
X_08342_ _09150_/A _11798_/A VGND VGND VPWR VPWR _08364_/A sky130_fd_sc_hd__or2_2
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08273_ _08307_/A VGND VGND VPWR VPWR _08292_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07224_ _07277_/B _07161_/B _07223_/X _07220_/Y VGND VGND VPWR VPWR _15647_/D sky130_fd_sc_hd__a211oi_1
X_07155_ _07285_/B _07233_/A VGND VGND VPWR VPWR _07231_/A sky130_fd_sc_hd__or2_1
XFILLER_118_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07988_ _07988_/A VGND VGND VPWR VPWR _07988_/X sky130_fd_sc_hd__buf_1
XFILLER_28_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09727_ _09737_/A VGND VGND VPWR VPWR _09727_/X sky130_fd_sc_hd__buf_1
XFILLER_86_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09658_ _15019_/Q _09641_/X _09657_/X _09645_/X VGND VGND VPWR VPWR _15019_/D sky130_fd_sc_hd__a22o_1
XFILLER_15_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08609_ _15283_/Q _08607_/X _08448_/X _08608_/X VGND VGND VPWR VPWR _15283_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _10349_/A VGND VGND VPWR VPWR _09589_/X sky130_fd_sc_hd__buf_1
XFILLER_31_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11628_/A VGND VGND VPWR VPWR _11620_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _11556_/A VGND VGND VPWR VPWR _11551_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10502_ _14801_/Q _10496_/X _10375_/X _10497_/X VGND VGND VPWR VPWR _14801_/D sky130_fd_sc_hd__a22o_1
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _14949_/Q _15045_/Q _15013_/Q _15077_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14270_/X sky130_fd_sc_hd__mux4_2
X_11482_ _11508_/A VGND VGND VPWR VPWR _11493_/A sky130_fd_sc_hd__buf_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ _13222_/X _13232_/X _15562_/Q VGND VGND VPWR VPWR _13221_/X sky130_fd_sc_hd__mux2_1
X_10433_ _10433_/A VGND VGND VPWR VPWR _10433_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13152_ _12817_/B _12995_/Y _13152_/S VGND VGND VPWR VPWR _13152_/X sky130_fd_sc_hd__mux2_1
X_10364_ _14836_/Q _10353_/X _10363_/X _10356_/X VGND VGND VPWR VPWR _14836_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12103_ _12103_/A VGND VGND VPWR VPWR _12346_/A sky130_fd_sc_hd__buf_1
XFILLER_152_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13083_ _12342_/X _15585_/Q _13090_/S VGND VGND VPWR VPWR _13083_/X sky130_fd_sc_hd__mux2_1
X_10295_ _10311_/A VGND VGND VPWR VPWR _10296_/A sky130_fd_sc_hd__buf_1
XFILLER_105_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12034_ _15520_/Q VGND VGND VPWR VPWR _12984_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13985_ _15137_/Q _15361_/Q _15329_/Q _15297_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13985_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12936_ _12765_/X _12763_/X _12919_/D _12935_/X VGND VGND VPWR VPWR _12937_/B sky130_fd_sc_hd__o22a_1
XFILLER_46_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12867_ _12867_/A _12867_/B VGND VGND VPWR VPWR _12867_/Y sky130_fd_sc_hd__nor2_1
X_15655_ _15669_/CLK _15655_/D VGND VGND VPWR VPWR _15655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14606_ _11278_/X _14606_/D VGND VGND VPWR VPWR _14606_/Q sky130_fd_sc_hd__dfxtp_1
X_11818_ _11818_/A VGND VGND VPWR VPWR _11818_/X sky130_fd_sc_hd__clkbuf_1
X_15586_ _15590_/CLK _15586_/D VGND VGND VPWR VPWR _15586_/Q sky130_fd_sc_hd__dfxtp_1
X_12798_ _12798_/A VGND VGND VPWR VPWR _12798_/X sky130_fd_sc_hd__buf_1
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14537_ _11544_/X _14537_/D VGND VGND VPWR VPWR _14537_/Q sky130_fd_sc_hd__dfxtp_1
X_11749_ _11751_/A VGND VGND VPWR VPWR _11749_/X sky130_fd_sc_hd__clkbuf_1
X_14468_ _11792_/X _14468_/D VGND VGND VPWR VPWR _14468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13419_ _12976_/Y _12963_/X _13419_/S VGND VGND VPWR VPWR _13419_/X sky130_fd_sc_hd__mux2_1
X_14399_ _14399_/CLK instruction[15] VGND VGND VPWR VPWR _14399_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08960_ _15194_/Q _08954_/X _08822_/X _08955_/X VGND VGND VPWR VPWR _15194_/D sky130_fd_sc_hd__a22o_1
XFILLER_142_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clkbuf_opt_3_clk/X VGND VGND VPWR VPWR _14401_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07911_ _07910_/A _07760_/B _07910_/Y _15593_/Q _07835_/X VGND VGND VPWR VPWR _15427_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_142_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08891_ _09263_/A VGND VGND VPWR VPWR _08891_/X sky130_fd_sc_hd__buf_1
X_07842_ _07813_/X _07683_/X _07841_/X VGND VGND VPWR VPWR _07843_/A sky130_fd_sc_hd__o21ai_1
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07773_ _07772_/A _07873_/A _07733_/Y _07734_/X _07772_/X VGND VGND VPWR VPWR _07856_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_84_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09512_ _15046_/Q _09505_/X _09279_/X _09506_/X VGND VGND VPWR VPWR _15046_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09443_ _15066_/Q _09436_/X _09192_/X _09437_/X VGND VGND VPWR VPWR _15066_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09374_ _09374_/A VGND VGND VPWR VPWR _09395_/A sky130_fd_sc_hd__clkbuf_2
X_08325_ _08325_/A VGND VGND VPWR VPWR _08325_/X sky130_fd_sc_hd__buf_1
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08256_ _08260_/A VGND VGND VPWR VPWR _08256_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07207_ _07265_/B _07169_/B _07200_/X _07205_/Y VGND VGND VPWR VPWR _15655_/D sky130_fd_sc_hd__a211oi_2
XFILLER_119_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08187_ _08189_/A VGND VGND VPWR VPWR _08187_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07138_ _13106_/X VGND VGND VPWR VPWR _07269_/B sky130_fd_sc_hd__inv_2
XFILLER_134_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10080_ _10173_/A VGND VGND VPWR VPWR _10143_/A sky130_fd_sc_hd__buf_1
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13770_ _14967_/Q _15063_/Q _15031_/Q _15095_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13770_/X sky130_fd_sc_hd__mux4_1
X_10982_ _10984_/A VGND VGND VPWR VPWR _10982_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12721_ _12735_/A _12735_/B VGND VGND VPWR VPWR _12721_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15440_ _15667_/CLK _15440_/D VGND VGND VPWR VPWR data_address[13] sky130_fd_sc_hd__dfxtp_4
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _12652_/A VGND VGND VPWR VPWR _12652_/X sky130_fd_sc_hd__buf_1
XFILLER_90_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _11612_/A VGND VGND VPWR VPWR _11603_/X sky130_fd_sc_hd__buf_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ _08189_/X _15371_/D VGND VGND VPWR VPWR _15371_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ _12579_/X _12625_/A _12625_/B _12286_/A VGND VGND VPWR VPWR _12598_/B sky130_fd_sc_hd__a31o_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14322_ _15505_/CLK _14322_/D VGND VGND VPWR VPWR _14322_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ _14540_/Q _11527_/X _11533_/X _11530_/X VGND VGND VPWR VPWR _14540_/D sky130_fd_sc_hd__a22o_1
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ _14662_/Q _15238_/Q _14726_/Q _14694_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14253_/X sky130_fd_sc_hd__mux4_2
X_11465_ _14556_/Q _11462_/X _11463_/X _11464_/X VGND VGND VPWR VPWR _14556_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13204_ _13203_/X _12824_/X _15565_/Q VGND VGND VPWR VPWR _13204_/X sky130_fd_sc_hd__mux2_1
X_10416_ _14824_/Q _10406_/X _10415_/X _10408_/X VGND VGND VPWR VPWR _14824_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14184_ _15181_/Q _15149_/Q _14765_/Q _14797_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14184_/X sky130_fd_sc_hd__mux4_1
X_11396_ _11415_/A VGND VGND VPWR VPWR _11396_/X sky130_fd_sc_hd__buf_1
XFILLER_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13135_ _12138_/X _13012_/Y _13152_/S VGND VGND VPWR VPWR _13135_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10347_ _10373_/A VGND VGND VPWR VPWR _10358_/A sky130_fd_sc_hd__buf_1
XFILLER_140_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13066_ _12814_/Y _15568_/Q _13076_/S VGND VGND VPWR VPWR _13066_/X sky130_fd_sc_hd__mux2_2
XFILLER_97_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10278_ _14856_/Q _10267_/X _10047_/X _10268_/X VGND VGND VPWR VPWR _14856_/D sky130_fd_sc_hd__a22o_1
X_12017_ _12017_/A VGND VGND VPWR VPWR _12017_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13968_ _14499_/Q _14467_/Q _14435_/Q _14403_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13968_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12919_ _12919_/A _12937_/A _12919_/C _12919_/D VGND VGND VPWR VPWR _12958_/A sky130_fd_sc_hd__or4_4
XFILLER_80_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13899_ _14826_/Q _14858_/Q _14890_/Q _14922_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13899_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15638_ _15669_/CLK _15638_/D VGND VGND VPWR VPWR _15638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15569_ _15578_/CLK _15569_/D VGND VGND VPWR VPWR _15569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08110_ _08120_/A VGND VGND VPWR VPWR _08123_/A sky130_fd_sc_hd__inv_2
X_09090_ _09094_/A VGND VGND VPWR VPWR _09090_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08041_ _14315_/Q VGND VGND VPWR VPWR _08042_/A sky130_fd_sc_hd__buf_1
XFILLER_147_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09992_ _14933_/Q _09985_/X _09991_/X _09988_/X VGND VGND VPWR VPWR _14933_/D sky130_fd_sc_hd__a22o_1
XFILLER_115_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08943_ _08963_/A VGND VGND VPWR VPWR _08943_/X sky130_fd_sc_hd__buf_1
X_08874_ _15214_/Q _08864_/X _08873_/X _08866_/X VGND VGND VPWR VPWR _15214_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07825_ _07813_/X _07688_/X _07831_/B VGND VGND VPWR VPWR _07826_/A sky130_fd_sc_hd__o21ai_1
XFILLER_57_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07756_ _07756_/A _15595_/Q VGND VGND VPWR VPWR _07756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07687_ _07687_/A _13132_/X VGND VGND VPWR VPWR _07695_/A sky130_fd_sc_hd__or2_2
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09426_ _09426_/A VGND VGND VPWR VPWR _09487_/A sky130_fd_sc_hd__buf_2
XFILLER_40_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09357_ _09366_/A VGND VGND VPWR VPWR _09357_/X sky130_fd_sc_hd__buf_1
XFILLER_100_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08308_ _08326_/A VGND VGND VPWR VPWR _08308_/X sky130_fd_sc_hd__buf_1
X_09288_ _15108_/Q _09152_/A _09287_/X _09156_/A VGND VGND VPWR VPWR _15108_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08239_ _08239_/A VGND VGND VPWR VPWR _08305_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_153_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11250_ _11310_/A VGND VGND VPWR VPWR _11271_/A sky130_fd_sc_hd__buf_2
XFILLER_119_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10201_ _10201_/A VGND VGND VPWR VPWR _10206_/A sky130_fd_sc_hd__buf_1
XFILLER_122_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11181_ _11203_/A VGND VGND VPWR VPWR _11190_/A sky130_fd_sc_hd__buf_1
XFILLER_107_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10132_ _10132_/A VGND VGND VPWR VPWR _10132_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10063_ _14916_/Q _09927_/A _10062_/X _09931_/A VGND VGND VPWR VPWR _14916_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14940_ _09956_/X _14940_/D VGND VGND VPWR VPWR _14940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14871_ _10223_/X _14871_/D VGND VGND VPWR VPWR _14871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13822_ _15217_/Q _14545_/Q _14993_/Q _15409_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13822_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13753_ _14680_/Q _15256_/Q _14744_/Q _14712_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13753_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10965_ _10965_/A VGND VGND VPWR VPWR _11026_/A sky130_fd_sc_hd__buf_4
XFILLER_141_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12704_ _13243_/X _12698_/X _13238_/X _12701_/X _12703_/X VGND VGND VPWR VPWR _12704_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_44_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13684_ _15199_/Q _15167_/Q _14783_/Q _14815_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13684_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10896_ _14707_/Q _10894_/X _10751_/X _10895_/X VGND VGND VPWR VPWR _14707_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ _12635_/A VGND VGND VPWR VPWR _12635_/X sky130_fd_sc_hd__clkbuf_4
X_15423_ _07946_/X _15423_/D VGND VGND VPWR VPWR _15423_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15354_ _08258_/X _15354_/D VGND VGND VPWR VPWR _15354_/Q sky130_fd_sc_hd__dfxtp_1
X_12566_ _12563_/C _12565_/X _07301_/X VGND VGND VPWR VPWR _12575_/B sky130_fd_sc_hd__o21a_1
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _11517_/A VGND VGND VPWR VPWR _11517_/X sky130_fd_sc_hd__clkbuf_1
X_14305_ _15521_/CLK _14305_/D VGND VGND VPWR VPWR _14305_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15285_ _08601_/X _15285_/D VGND VGND VPWR VPWR _15285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12497_ _12951_/A _12492_/X _12336_/X _12496_/X _12489_/X VGND VGND VPWR VPWR _12497_/X
+ sky130_fd_sc_hd__o32a_1
X_14236_ _14232_/X _14233_/X _14234_/X _14235_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14236_/X sky130_fd_sc_hd__mux4_2
X_11448_ _11474_/A VGND VGND VPWR VPWR _11448_/X sky130_fd_sc_hd__buf_1
XFILLER_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14167_ _14639_/Q _14607_/Q _14575_/Q _15375_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14167_/X sky130_fd_sc_hd__mux4_2
X_11379_ _11383_/A VGND VGND VPWR VPWR _11379_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13118_ _15664_/Q data_address[29] _15667_/Q VGND VGND VPWR VPWR _13118_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14098_ _14518_/Q _14486_/Q _14454_/Q _14422_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14098_/X sky130_fd_sc_hd__mux4_1
X_13049_ wdata[22] rdata[22] _13057_/S VGND VGND VPWR VPWR _14326_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07610_ _07638_/A _13061_/X VGND VGND VPWR VPWR _15476_/D sky130_fd_sc_hd__and2_1
X_08590_ _08592_/A VGND VGND VPWR VPWR _08590_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07541_ _07541_/A VGND VGND VPWR VPWR _07541_/Y sky130_fd_sc_hd__inv_2
X_07472_ _07472_/A _13490_/X VGND VGND VPWR VPWR _15540_/D sky130_fd_sc_hd__and2_1
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09211_ _09211_/A VGND VGND VPWR VPWR _09211_/X sky130_fd_sc_hd__buf_1
X_09142_ _09144_/A VGND VGND VPWR VPWR _09142_/X sky130_fd_sc_hd__clkbuf_1
X_09073_ _15162_/Q _09065_/X _08822_/X _09066_/X VGND VGND VPWR VPWR _15162_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08024_ _08034_/A VGND VGND VPWR VPWR _08024_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09975_ _14937_/Q _09972_/X _09973_/X _09974_/X VGND VGND VPWR VPWR _14937_/D sky130_fd_sc_hd__a22o_1
XFILLER_131_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08926_ _10548_/B VGND VGND VPWR VPWR _10438_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_130_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08857_ _15218_/Q _08851_/X _08856_/X _08853_/X VGND VGND VPWR VPWR _15218_/D sky130_fd_sc_hd__a22o_1
XFILLER_73_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07808_ _07808_/A VGND VGND VPWR VPWR _07808_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08788_ _08788_/A VGND VGND VPWR VPWR _08788_/X sky130_fd_sc_hd__clkbuf_1
X_07739_ _07769_/A VGND VGND VPWR VPWR _07739_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10750_ _10750_/A VGND VGND VPWR VPWR _11502_/A sky130_fd_sc_hd__buf_2
XFILLER_53_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09409_ _09423_/A VGND VGND VPWR VPWR _09410_/A sky130_fd_sc_hd__buf_1
X_10681_ _10779_/A VGND VGND VPWR VPWR _10716_/A sky130_fd_sc_hd__clkbuf_2
X_12420_ _12904_/D VGND VGND VPWR VPWR _12420_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12351_ _12355_/A VGND VGND VPWR VPWR _12363_/A sky130_fd_sc_hd__buf_1
XFILLER_138_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11302_ _11308_/A VGND VGND VPWR VPWR _11302_/X sky130_fd_sc_hd__clkbuf_1
X_15070_ _09431_/X _15070_/D VGND VGND VPWR VPWR _15070_/Q sky130_fd_sc_hd__dfxtp_1
X_12282_ _12162_/Y _12273_/Y _12177_/Y _12279_/X _12281_/X VGND VGND VPWR VPWR _12282_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14021_ _14017_/X _14018_/X _14019_/X _14020_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14021_/X sky130_fd_sc_hd__mux4_1
X_11233_ _11242_/A VGND VGND VPWR VPWR _11233_/X sky130_fd_sc_hd__buf_1
XFILLER_136_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11164_ _14637_/Q _11160_/X _11161_/X _11163_/X VGND VGND VPWR VPWR _14637_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10115_ _10123_/A VGND VGND VPWR VPWR _10115_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11095_ _11463_/A VGND VGND VPWR VPWR _11095_/X sky130_fd_sc_hd__buf_1
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14923_ _10033_/X _14923_/D VGND VGND VPWR VPWR _14923_/Q sky130_fd_sc_hd__dfxtp_1
X_10046_ _10054_/A VGND VGND VPWR VPWR _10046_/X sky130_fd_sc_hd__buf_1
XFILLER_76_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14854_ _10284_/X _14854_/D VGND VGND VPWR VPWR _14854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13805_ _15123_/Q _15347_/Q _15315_/Q _15283_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13805_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11997_ _12006_/A VGND VGND VPWR VPWR _11997_/X sky130_fd_sc_hd__buf_1
X_14785_ _10557_/X _14785_/D VGND VGND VPWR VPWR _14785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10948_ _10948_/A VGND VGND VPWR VPWR _10948_/X sky130_fd_sc_hd__clkbuf_1
X_13736_ _13732_/X _13733_/X _13734_/X _13735_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13736_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10879_ _10879_/A VGND VGND VPWR VPWR _10879_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13667_ _14657_/Q _14625_/Q _14593_/Q _15393_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13667_/X sky130_fd_sc_hd__mux4_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15406_ _08040_/X _15406_/D VGND VGND VPWR VPWR _15406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12618_ _12618_/A VGND VGND VPWR VPWR _12618_/X sky130_fd_sc_hd__buf_1
X_13598_ _13597_/X _14317_/D _15506_/Q VGND VGND VPWR VPWR _13598_/X sky130_fd_sc_hd__mux2_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12549_ _12556_/A _12559_/B VGND VGND VPWR VPWR _12549_/Y sky130_fd_sc_hd__nor2_1
X_15337_ _08320_/X _15337_/D VGND VGND VPWR VPWR _15337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 data_address[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15268_ _08655_/X _15268_/D VGND VGND VPWR VPWR _15268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14219_ _14826_/Q _14858_/Q _14890_/Q _14922_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14219_/X sky130_fd_sc_hd__mux4_2
X_15199_ _08940_/X _15199_/D VGND VGND VPWR VPWR _15199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09760_ _14994_/Q _09756_/X _09617_/X _09757_/X VGND VGND VPWR VPWR _14994_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08711_ _08741_/A VGND VGND VPWR VPWR _08732_/A sky130_fd_sc_hd__buf_1
X_09691_ _10431_/A VGND VGND VPWR VPWR _09691_/X sky130_fd_sc_hd__buf_1
XFILLER_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08642_ _08642_/A VGND VGND VPWR VPWR _08642_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08573_ _15293_/Q _08565_/X _08384_/X _08568_/X VGND VGND VPWR VPWR _15293_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07524_ _07524_/A VGND VGND VPWR VPWR _11559_/A sky130_fd_sc_hd__buf_1
XFILLER_23_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07455_ _07455_/A _13454_/X VGND VGND VPWR VPWR _15552_/D sky130_fd_sc_hd__and2_1
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07386_ _13157_/X VGND VGND VPWR VPWR _07386_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09125_ _09125_/A VGND VGND VPWR VPWR _09125_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09056_ _09117_/A VGND VGND VPWR VPWR _09076_/A sky130_fd_sc_hd__clkbuf_2
X_08007_ _15413_/Q _07998_/X _08006_/X _08002_/X VGND VGND VPWR VPWR _15413_/D sky130_fd_sc_hd__a22o_1
XFILLER_151_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09958_ _10328_/A VGND VGND VPWR VPWR _09958_/X sky130_fd_sc_hd__buf_1
XFILLER_58_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08909_ _09279_/A VGND VGND VPWR VPWR _08909_/X sky130_fd_sc_hd__buf_1
XFILLER_46_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09889_ _09908_/A VGND VGND VPWR VPWR _09889_/X sky130_fd_sc_hd__buf_1
XFILLER_57_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11920_ _14432_/Q _11912_/X _07944_/A _11915_/X VGND VGND VPWR VPWR _14432_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11851_ _11907_/A VGND VGND VPWR VPWR _11870_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_122_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10802_ _10802_/A VGND VGND VPWR VPWR _10802_/X sky130_fd_sc_hd__clkbuf_1
X_14570_ _11403_/X _14570_/D VGND VGND VPWR VPWR _14570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11782_ _11782_/A VGND VGND VPWR VPWR _11782_/X sky130_fd_sc_hd__clkbuf_1
X_13521_ _13966_/X _13971_/X _13521_/S VGND VGND VPWR VPWR _13521_/X sky130_fd_sc_hd__mux2_1
X_10733_ _10733_/A VGND VGND VPWR VPWR _11489_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13452_ _13736_/X _13741_/X _14386_/Q VGND VGND VPWR VPWR _13452_/X sky130_fd_sc_hd__mux2_2
X_10664_ _10664_/A VGND VGND VPWR VPWR _11431_/A sky130_fd_sc_hd__buf_1
X_12403_ _15588_/Q VGND VGND VPWR VPWR _12403_/X sky130_fd_sc_hd__buf_1
X_13383_ _12812_/A _12775_/X _13418_/S VGND VGND VPWR VPWR _13383_/X sky130_fd_sc_hd__mux2_1
X_10595_ _10595_/A VGND VGND VPWR VPWR _10595_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12334_ _12478_/A VGND VGND VPWR VPWR _12739_/A sky130_fd_sc_hd__buf_1
X_15122_ _09227_/X _15122_/D VGND VGND VPWR VPWR _15122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15053_ _09484_/X _15053_/D VGND VGND VPWR VPWR _15053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12265_ _12265_/A VGND VGND VPWR VPWR _12802_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14004_ _15199_/Q _15167_/Q _14783_/Q _14815_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14004_/X sky130_fd_sc_hd__mux4_2
X_11216_ _11216_/A VGND VGND VPWR VPWR _11239_/A sky130_fd_sc_hd__buf_2
XFILLER_141_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12196_ _15569_/Q VGND VGND VPWR VPWR _12788_/A sky130_fd_sc_hd__inv_2
X_11147_ _11147_/A VGND VGND VPWR VPWR _11147_/X sky130_fd_sc_hd__buf_1
XFILLER_68_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11078_ _11078_/A VGND VGND VPWR VPWR _11159_/A sky130_fd_sc_hd__buf_2
XFILLER_83_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10029_ _10029_/A VGND VGND VPWR VPWR _10029_/X sky130_fd_sc_hd__clkbuf_1
X_14906_ _10102_/X _14906_/D VGND VGND VPWR VPWR _14906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14837_ _10358_/X _14837_/D VGND VGND VPWR VPWR _14837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14768_ _10615_/X _14768_/D VGND VGND VPWR VPWR _14768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13719_ _14844_/Q _14876_/Q _14908_/Q _14940_/Q _13740_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13719_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14699_ _10920_/X _14699_/D VGND VGND VPWR VPWR _14699_/Q sky130_fd_sc_hd__dfxtp_1
X_07240_ _07240_/A VGND VGND VPWR VPWR _07288_/B sky130_fd_sc_hd__buf_1
XFILLER_118_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07171_ _07263_/B _07171_/B VGND VGND VPWR VPWR _07202_/A sky130_fd_sc_hd__or2_1
XFILLER_118_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09812_ _09812_/A VGND VGND VPWR VPWR _09812_/X sky130_fd_sc_hd__buf_1
XFILLER_86_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09743_ _09754_/A VGND VGND VPWR VPWR _09752_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09674_ _09680_/A VGND VGND VPWR VPWR _09674_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08625_ _08633_/A VGND VGND VPWR VPWR _08625_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08556_ _15298_/Q _08552_/X _08347_/X _08555_/X VGND VGND VPWR VPWR _15298_/D sky130_fd_sc_hd__a22o_1
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07507_ _07511_/A VGND VGND VPWR VPWR _07510_/A sky130_fd_sc_hd__buf_1
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08487_ _08524_/A VGND VGND VPWR VPWR _08487_/X sky130_fd_sc_hd__buf_1
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07438_ _07438_/A _13639_/X VGND VGND VPWR VPWR _15564_/D sky130_fd_sc_hd__and2_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07369_ _07370_/B VGND VGND VPWR VPWR _07369_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09108_ _15152_/Q _09106_/X _08865_/X _09107_/X VGND VGND VPWR VPWR _15152_/D sky130_fd_sc_hd__a22o_1
X_10380_ _10380_/A VGND VGND VPWR VPWR _10380_/X sky130_fd_sc_hd__buf_1
XFILLER_108_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09039_ _09408_/A _10438_/B VGND VGND VPWR VPWR _09052_/A sky130_fd_sc_hd__or2_2
X_12050_ _12977_/A _12050_/B VGND VGND VPWR VPWR _13425_/S sky130_fd_sc_hd__nor2_4
XFILLER_77_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11001_ _11005_/A VGND VGND VPWR VPWR _11001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12952_ _12905_/A _12903_/X _12959_/C _12950_/X _12951_/X VGND VGND VPWR VPWR _12952_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_133_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11903_ _11905_/A VGND VGND VPWR VPWR _11903_/X sky130_fd_sc_hd__clkbuf_1
X_15671_ _15672_/D _12992_/Y VGND VGND VPWR VPWR _15671_/Q sky130_fd_sc_hd__dlxtn_1
X_12883_ _12883_/A _12883_/B VGND VGND VPWR VPWR _12884_/A sky130_fd_sc_hd__or2_1
XANTENNA_210 _13498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_221 _15453_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_232 _09577_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_243 _11587_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14622_ _11226_/X _14622_/D VGND VGND VPWR VPWR _14622_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_254 _12745_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11834_ _11834_/A VGND VGND VPWR VPWR _11834_/X sky130_fd_sc_hd__buf_1
XFILLER_14_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11765_ _11765_/A VGND VGND VPWR VPWR _11784_/A sky130_fd_sc_hd__buf_1
X_14553_ _11473_/X _14553_/D VGND VGND VPWR VPWR _14553_/Q sky130_fd_sc_hd__dfxtp_1
X_10716_ _10716_/A VGND VGND VPWR VPWR _10716_/X sky130_fd_sc_hd__buf_1
X_13504_ _13503_/X rdata[6] _13516_/S VGND VGND VPWR VPWR _13504_/X sky130_fd_sc_hd__mux2_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14484_ _11740_/X _14484_/D VGND VGND VPWR VPWR _14484_/Q sky130_fd_sc_hd__dfxtp_1
X_11696_ _14497_/Q _11688_/X _11437_/X _11691_/X VGND VGND VPWR VPWR _14497_/D sky130_fd_sc_hd__a22o_1
X_13435_ _13434_/X rdata[29] _13516_/S VGND VGND VPWR VPWR _13435_/X sky130_fd_sc_hd__mux2_1
X_10647_ _10647_/A VGND VGND VPWR VPWR _10647_/X sky130_fd_sc_hd__buf_1
XFILLER_10_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13366_ _12415_/X _12435_/X _13418_/S VGND VGND VPWR VPWR _13366_/X sky130_fd_sc_hd__mux2_1
X_10578_ _10578_/A VGND VGND VPWR VPWR _10583_/A sky130_fd_sc_hd__buf_1
X_15105_ _09303_/X _15105_/D VGND VGND VPWR VPWR _15105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12317_ _12699_/A _12740_/A VGND VGND VPWR VPWR _12367_/A sky130_fd_sc_hd__or2_1
X_13297_ _12820_/X _12847_/A _13418_/S VGND VGND VPWR VPWR _13297_/X sky130_fd_sc_hd__mux2_1
X_12248_ _12820_/A _12246_/B _12247_/Y VGND VGND VPWR VPWR _12265_/A sky130_fd_sc_hd__a21oi_1
X_15036_ _09561_/X _15036_/D VGND VGND VPWR VPWR _15036_/Q sky130_fd_sc_hd__dfxtp_1
X_12179_ _15572_/Q VGND VGND VPWR VPWR _12179_/X sky130_fd_sc_hd__buf_1
XFILLER_68_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08410_ _15321_/Q _08405_/X _08408_/X _08409_/X VGND VGND VPWR VPWR _15321_/D sky130_fd_sc_hd__a22o_1
X_09390_ _15081_/Q _09386_/X _09267_/X _09387_/X VGND VGND VPWR VPWR _15081_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08341_ _09521_/A VGND VGND VPWR VPWR _11798_/A sky130_fd_sc_hd__buf_1
XFILLER_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08272_ _08291_/A VGND VGND VPWR VPWR _08272_/X sky130_fd_sc_hd__buf_1
XFILLER_149_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07223_ _07246_/A VGND VGND VPWR VPWR _07223_/X sky130_fd_sc_hd__buf_1
XFILLER_149_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07154_ _07236_/A _07237_/A _07242_/A _07286_/B VGND VGND VPWR VPWR _07233_/A sky130_fd_sc_hd__or4_4
XFILLER_146_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07987_ _14325_/Q VGND VGND VPWR VPWR _07988_/A sky130_fd_sc_hd__buf_1
XFILLER_47_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09726_ _09736_/A VGND VGND VPWR VPWR _09726_/X sky130_fd_sc_hd__buf_1
XFILLER_28_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09657_ _10403_/A VGND VGND VPWR VPWR _09657_/X sky130_fd_sc_hd__buf_1
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08608_ _08618_/A VGND VGND VPWR VPWR _08608_/X sky130_fd_sc_hd__buf_1
X_09588_ _10727_/A VGND VGND VPWR VPWR _10349_/A sky130_fd_sc_hd__buf_1
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _10827_/A VGND VGND VPWR VPWR _09287_/A sky130_fd_sc_hd__buf_1
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _14536_/Q _11540_/X _11549_/X _11542_/X VGND VGND VPWR VPWR _14536_/D sky130_fd_sc_hd__a22o_1
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10501_ _10501_/A VGND VGND VPWR VPWR _10501_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11481_ _11520_/A VGND VGND VPWR VPWR _11508_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ _13221_/X _13240_/X _13408_/S VGND VGND VPWR VPWR _13220_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10432_ _14820_/Q _10296_/A _10431_/X _10300_/A VGND VGND VPWR VPWR _14820_/D sky130_fd_sc_hd__a22o_1
XFILLER_109_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13151_ _12885_/X _12996_/Y _13152_/S VGND VGND VPWR VPWR _13151_/X sky130_fd_sc_hd__mux2_1
X_10363_ _10363_/A VGND VGND VPWR VPWR _10363_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_152_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12102_ _12102_/A VGND VGND VPWR VPWR _12103_/A sky130_fd_sc_hd__buf_1
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13082_ _12597_/Y _15584_/Q _13090_/S VGND VGND VPWR VPWR _13082_/X sky130_fd_sc_hd__mux2_1
X_10294_ _10294_/A _10294_/B VGND VGND VPWR VPWR _10311_/A sky130_fd_sc_hd__or2_1
XFILLER_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12033_ _12337_/A VGND VGND VPWR VPWR _12316_/A sky130_fd_sc_hd__inv_2
XFILLER_88_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13984_ _15201_/Q _15169_/Q _14785_/Q _14817_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13984_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12935_ _12791_/X _12788_/A _12919_/A _12778_/X _12785_/B VGND VGND VPWR VPWR _12935_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_34_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15654_ _15654_/CLK _15654_/D VGND VGND VPWR VPWR _15654_/Q sky130_fd_sc_hd__dfxtp_1
X_12866_ _15532_/Q VGND VGND VPWR VPWR _12867_/B sky130_fd_sc_hd__buf_1
XFILLER_34_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14605_ _11282_/X _14605_/D VGND VGND VPWR VPWR _14605_/Q sky130_fd_sc_hd__dfxtp_1
X_11817_ _14463_/Q _11813_/X _07951_/A _11816_/X VGND VGND VPWR VPWR _14463_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15585_ _15590_/CLK _15585_/D VGND VGND VPWR VPWR _15585_/Q sky130_fd_sc_hd__dfxtp_1
X_12797_ _12929_/A _12797_/B VGND VGND VPWR VPWR _12883_/B sky130_fd_sc_hd__nand2_1
XFILLER_42_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14536_ _11548_/X _14536_/D VGND VGND VPWR VPWR _14536_/Q sky130_fd_sc_hd__dfxtp_1
X_11748_ _14482_/Q _11743_/X _11506_/X _11744_/X VGND VGND VPWR VPWR _14482_/D sky130_fd_sc_hd__a22o_1
XFILLER_41_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14467_ _11795_/X _14467_/D VGND VGND VPWR VPWR _14467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11679_ _14501_/Q _11673_/X _11564_/X _11674_/X VGND VGND VPWR VPWR _14501_/D sky130_fd_sc_hd__a22o_1
XFILLER_146_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13418_ _12875_/B _12211_/X _13418_/S VGND VGND VPWR VPWR _13418_/X sky130_fd_sc_hd__mux2_1
X_14398_ _15652_/CLK instruction[23] VGND VGND VPWR VPWR _14398_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13349_ _13406_/X _13404_/X _13415_/S VGND VGND VPWR VPWR _13349_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07910_ _07910_/A VGND VGND VPWR VPWR _07910_/Y sky130_fd_sc_hd__inv_2
X_15019_ _09655_/X _15019_/D VGND VGND VPWR VPWR _15019_/Q sky130_fd_sc_hd__dfxtp_1
X_08890_ _08904_/A VGND VGND VPWR VPWR _08890_/X sky130_fd_sc_hd__buf_1
X_07841_ _07841_/A _07846_/A VGND VGND VPWR VPWR _07841_/X sky130_fd_sc_hd__or2_1
XFILLER_69_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07772_ _07772_/A _07873_/A _07772_/C _07876_/A VGND VGND VPWR VPWR _07772_/X sky130_fd_sc_hd__or4b_4
XFILLER_83_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09511_ _09515_/A VGND VGND VPWR VPWR _09511_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09442_ _09444_/A VGND VGND VPWR VPWR _09442_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09373_ _09381_/A VGND VGND VPWR VPWR _09373_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08324_ _08324_/A VGND VGND VPWR VPWR _08324_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08255_ _08255_/A VGND VGND VPWR VPWR _08260_/A sky130_fd_sc_hd__buf_1
XFILLER_138_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07206_ _13110_/X _07205_/Y _07198_/X _07171_/B VGND VGND VPWR VPWR _15656_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08186_ _15373_/Q _08183_/X _08048_/X _08185_/X VGND VGND VPWR VPWR _15373_/D sky130_fd_sc_hd__a22o_1
XFILLER_118_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07137_ _13107_/X VGND VGND VPWR VPWR _07268_/B sky130_fd_sc_hd__inv_2
XFILLER_106_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09709_ _09709_/A VGND VGND VPWR VPWR _09709_/X sky130_fd_sc_hd__clkbuf_1
X_10981_ _14683_/Q _10976_/X _10708_/X _10977_/X VGND VGND VPWR VPWR _14683_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12720_ _12720_/A VGND VGND VPWR VPWR _12737_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12651_ _12651_/A _12651_/B VGND VGND VPWR VPWR _12651_/Y sky130_fd_sc_hd__nor2_1
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _11608_/A VGND VGND VPWR VPWR _11602_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ _12581_/X _12144_/X _12292_/X VGND VGND VPWR VPWR _12625_/B sky130_fd_sc_hd__o21ai_1
X_15370_ _08194_/X _15370_/D VGND VGND VPWR VPWR _15370_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14321_ _15517_/CLK _14321_/D VGND VGND VPWR VPWR _14321_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _11533_/A VGND VGND VPWR VPWR _11533_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14252_ _15206_/Q _14534_/Q _14982_/Q _15398_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14252_/X sky130_fd_sc_hd__mux4_2
X_11464_ _11476_/A VGND VGND VPWR VPWR _11464_/X sky130_fd_sc_hd__buf_1
XFILLER_137_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13203_ _13205_/X _13245_/X _13393_/S VGND VGND VPWR VPWR _13203_/X sky130_fd_sc_hd__mux2_1
X_10415_ _10415_/A VGND VGND VPWR VPWR _10415_/X sky130_fd_sc_hd__buf_1
X_14183_ _14669_/Q _15245_/Q _14733_/Q _14701_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14183_/X sky130_fd_sc_hd__mux4_2
X_11395_ _11395_/A VGND VGND VPWR VPWR _11415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13134_ _12635_/X _13013_/Y _13152_/S VGND VGND VPWR VPWR _13134_/X sky130_fd_sc_hd__mux2_1
X_10346_ _10346_/A VGND VGND VPWR VPWR _10373_/A sky130_fd_sc_hd__buf_2
XFILLER_125_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13065_ _12834_/Y _15567_/Q _13076_/S VGND VGND VPWR VPWR _13065_/X sky130_fd_sc_hd__mux2_2
X_10277_ _10279_/A VGND VGND VPWR VPWR _10277_/X sky130_fd_sc_hd__clkbuf_1
X_12016_ _14403_/Q _11912_/A _08099_/A _11915_/A VGND VGND VPWR VPWR _14403_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13967_ _14627_/Q _14595_/Q _14563_/Q _15363_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13967_/X sky130_fd_sc_hd__mux4_1
XFILLER_81_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12918_ _12765_/X _12187_/X _12762_/A _12763_/A VGND VGND VPWR VPWR _12919_/D sky130_fd_sc_hd__o22a_1
XFILLER_46_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13898_ _14506_/Q _14474_/Q _14442_/Q _14410_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13898_/X sky130_fd_sc_hd__mux4_2
X_15637_ _15648_/CLK _15637_/D VGND VGND VPWR VPWR _15637_/Q sky130_fd_sc_hd__dfxtp_1
X_12849_ _12349_/X _12841_/Y _12845_/Y _12848_/X VGND VGND VPWR VPWR _12849_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_15_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15568_ _15578_/CLK _15568_/D VGND VGND VPWR VPWR _15568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14519_ _11617_/X _14519_/D VGND VGND VPWR VPWR _14519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15499_ _15502_/CLK _15499_/D VGND VGND VPWR VPWR wdata[25] sky130_fd_sc_hd__dfxtp_1
X_08040_ _08052_/A VGND VGND VPWR VPWR _08040_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09991_ _10359_/A VGND VGND VPWR VPWR _09991_/X sky130_fd_sc_hd__buf_1
XFILLER_142_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08942_ _09005_/A VGND VGND VPWR VPWR _08963_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08873_ _09245_/A VGND VGND VPWR VPWR _08873_/X sky130_fd_sc_hd__buf_1
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07824_ _07830_/A _07830_/B VGND VGND VPWR VPWR _07831_/B sky130_fd_sc_hd__or2_1
XFILLER_111_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07755_ _13150_/X VGND VGND VPWR VPWR _07756_/A sky130_fd_sc_hd__inv_2
XFILLER_53_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07686_ _13131_/X VGND VGND VPWR VPWR _07686_/X sky130_fd_sc_hd__buf_1
XFILLER_25_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09425_ _09445_/A VGND VGND VPWR VPWR _09425_/X sky130_fd_sc_hd__buf_1
XFILLER_25_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09356_ _09365_/A VGND VGND VPWR VPWR _09356_/X sky130_fd_sc_hd__buf_1
X_08307_ _08307_/A VGND VGND VPWR VPWR _08326_/A sky130_fd_sc_hd__buf_1
X_09287_ _09287_/A VGND VGND VPWR VPWR _09287_/X sky130_fd_sc_hd__buf_1
XFILLER_100_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08238_ _08238_/A VGND VGND VPWR VPWR _08238_/X sky130_fd_sc_hd__buf_1
XFILLER_119_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08169_ _08169_/A VGND VGND VPWR VPWR _08169_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10200_ _14879_/Q _10196_/X _09944_/X _10199_/X VGND VGND VPWR VPWR _14879_/D sky130_fd_sc_hd__a22o_1
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11180_ _11216_/A VGND VGND VPWR VPWR _11203_/A sky130_fd_sc_hd__clkbuf_2
X_10131_ _14898_/Q _10127_/X _10003_/X _10128_/X VGND VGND VPWR VPWR _14898_/D sky130_fd_sc_hd__a22o_1
XFILLER_106_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10062_ _10431_/A VGND VGND VPWR VPWR _10062_/X sky130_fd_sc_hd__buf_1
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14870_ _10225_/X _14870_/D VGND VGND VPWR VPWR _14870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13821_ _13817_/X _13818_/X _13819_/X _13820_/X _07533_/A _13946_/S1 VGND VGND VPWR
+ VPWR _13821_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13752_ _15224_/Q _14552_/Q _15000_/Q _15416_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13752_/X sky130_fd_sc_hd__mux4_1
X_10964_ _10985_/A VGND VGND VPWR VPWR _10964_/X sky130_fd_sc_hd__buf_1
XFILLER_90_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12703_ _12703_/A _12703_/B _12758_/C VGND VGND VPWR VPWR _12703_/X sky130_fd_sc_hd__or3_2
X_13683_ _14687_/Q _15263_/Q _14751_/Q _14719_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13683_/X sky130_fd_sc_hd__mux4_2
X_10895_ _10905_/A VGND VGND VPWR VPWR _10895_/X sky130_fd_sc_hd__buf_1
X_15422_ _07956_/X _15422_/D VGND VGND VPWR VPWR _15422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ _12634_/A VGND VGND VPWR VPWR _12634_/X sky130_fd_sc_hd__clkbuf_4
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15353_ _08260_/X _15353_/D VGND VGND VPWR VPWR _15353_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12565_ _14394_/Q _14392_/Q _12565_/C VGND VGND VPWR VPWR _12565_/X sky130_fd_sc_hd__or3_4
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14304_ _15505_/CLK _14304_/D VGND VGND VPWR VPWR _14304_/Q sky130_fd_sc_hd__dfxtp_1
X_11516_ _14544_/Q _11513_/X _11514_/X _11515_/X VGND VGND VPWR VPWR _14544_/D sky130_fd_sc_hd__a22o_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15284_ _08603_/X _15284_/D VGND VGND VPWR VPWR _15284_/Q sky130_fd_sc_hd__dfxtp_1
X_12496_ _12620_/A VGND VGND VPWR VPWR _12496_/X sky130_fd_sc_hd__buf_1
XFILLER_8_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14235_ _15112_/Q _15336_/Q _15304_/Q _15272_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14235_/X sky130_fd_sc_hd__mux4_1
X_11447_ _11526_/A VGND VGND VPWR VPWR _11474_/A sky130_fd_sc_hd__clkbuf_2
X_11378_ _11398_/A VGND VGND VPWR VPWR _11383_/A sky130_fd_sc_hd__buf_1
X_14166_ _14162_/X _14163_/X _14164_/X _14165_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14166_/X sky130_fd_sc_hd__mux4_2
XFILLER_98_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13117_ _15663_/Q data_address[28] _15667_/Q VGND VGND VPWR VPWR _13117_/X sky130_fd_sc_hd__mux2_1
X_10329_ _10341_/A VGND VGND VPWR VPWR _10329_/X sky130_fd_sc_hd__buf_1
X_14097_ _14646_/Q _14614_/Q _14582_/Q _15382_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14097_/X sky130_fd_sc_hd__mux4_2
XFILLER_79_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13048_ wdata[21] rdata[21] _13057_/S VGND VGND VPWR VPWR _14325_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14999_ _09741_/X _14999_/D VGND VGND VPWR VPWR _14999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07540_ _15469_/Q VGND VGND VPWR VPWR _07540_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07471_ _07472_/A _13487_/X VGND VGND VPWR VPWR _15541_/D sky130_fd_sc_hd__and2_1
XFILLER_22_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09210_ _09235_/A VGND VGND VPWR VPWR _09210_/X sky130_fd_sc_hd__buf_1
X_09141_ _15142_/Q _09136_/X _08909_/X _09137_/X VGND VGND VPWR VPWR _15142_/D sky130_fd_sc_hd__a22o_1
XFILLER_147_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09072_ _09074_/A VGND VGND VPWR VPWR _09072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08023_ _08023_/A VGND VGND VPWR VPWR _08034_/A sky130_fd_sc_hd__buf_1
XFILLER_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09974_ _09974_/A VGND VGND VPWR VPWR _09974_/X sky130_fd_sc_hd__buf_1
XFILLER_130_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08925_ _08925_/A _09294_/B _08925_/C VGND VGND VPWR VPWR _10548_/B sky130_fd_sc_hd__or3_1
X_08856_ _09228_/A VGND VGND VPWR VPWR _08856_/X sky130_fd_sc_hd__buf_1
XFILLER_29_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07807_ _07807_/A VGND VGND VPWR VPWR _07807_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08787_ _15234_/Q _08782_/X _08783_/X _08786_/X VGND VGND VPWR VPWR _15234_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07738_ _13145_/X VGND VGND VPWR VPWR _07769_/A sky130_fd_sc_hd__inv_2
XFILLER_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07669_ _07675_/A VGND VGND VPWR VPWR _07781_/A sky130_fd_sc_hd__clkbuf_1
X_09408_ _09408_/A _09523_/B VGND VGND VPWR VPWR _09423_/A sky130_fd_sc_hd__or2_1
XFILLER_13_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10680_ _10680_/A VGND VGND VPWR VPWR _10779_/A sky130_fd_sc_hd__buf_4
X_09339_ _15096_/Q _09335_/X _09200_/X _09336_/X VGND VGND VPWR VPWR _15096_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12350_ _15554_/Q VGND VGND VPWR VPWR _12355_/A sky130_fd_sc_hd__inv_2
XFILLER_126_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11301_ _11301_/A VGND VGND VPWR VPWR _11308_/A sky130_fd_sc_hd__buf_1
X_12281_ _12693_/A _12150_/A _12151_/Y _12690_/A VGND VGND VPWR VPWR _12281_/X sky130_fd_sc_hd__o22a_1
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14020_ _14974_/Q _15070_/Q _15038_/Q _15102_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14020_/X sky130_fd_sc_hd__mux4_2
X_11232_ _11241_/A VGND VGND VPWR VPWR _11232_/X sky130_fd_sc_hd__buf_1
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11163_ _11188_/A VGND VGND VPWR VPWR _11163_/X sky130_fd_sc_hd__buf_1
XFILLER_134_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10114_ _10134_/A VGND VGND VPWR VPWR _10123_/A sky130_fd_sc_hd__buf_1
XFILLER_121_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11094_ _11107_/A VGND VGND VPWR VPWR _11094_/X sky130_fd_sc_hd__buf_1
XFILLER_76_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10045_ _10067_/A VGND VGND VPWR VPWR _10054_/A sky130_fd_sc_hd__buf_1
X_14922_ _10036_/X _14922_/D VGND VGND VPWR VPWR _14922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14853_ _10286_/X _14853_/D VGND VGND VPWR VPWR _14853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13804_ _15187_/Q _15155_/Q _14771_/Q _14803_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13804_/X sky130_fd_sc_hd__mux4_1
XFILLER_63_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14784_ _10559_/X _14784_/D VGND VGND VPWR VPWR _14784_/Q sky130_fd_sc_hd__dfxtp_1
X_11996_ _12005_/A VGND VGND VPWR VPWR _11996_/X sky130_fd_sc_hd__buf_1
XFILLER_44_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13735_ _15130_/Q _15354_/Q _15322_/Q _15290_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13735_/X sky130_fd_sc_hd__mux4_1
X_10947_ _14691_/Q _10840_/A _10832_/X _10843_/A VGND VGND VPWR VPWR _14691_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13666_ _13662_/X _13663_/X _13664_/X _13665_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13666_/X sky130_fd_sc_hd__mux4_2
X_10878_ _14712_/Q _10874_/X _10723_/X _10875_/X VGND VGND VPWR VPWR _14712_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15405_ _08044_/X _15405_/D VGND VGND VPWR VPWR _15405_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ _12615_/X _12101_/X _12616_/X VGND VGND VPWR VPWR _12617_/Y sky130_fd_sc_hd__o21ai_2
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ _13596_/X _07310_/Y _13649_/S VGND VGND VPWR VPWR _13597_/X sky130_fd_sc_hd__mux2_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15336_ _08322_/X _15336_/D VGND VGND VPWR VPWR _15336_/Q sky130_fd_sc_hd__dfxtp_1
X_12548_ _12545_/A _12551_/A data_address[0] VGND VGND VPWR VPWR _12559_/B sky130_fd_sc_hd__o21a_1
XFILLER_117_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15267_ _08657_/X _15267_/D VGND VGND VPWR VPWR _15267_/Q sky130_fd_sc_hd__dfxtp_1
X_12479_ _12784_/A VGND VGND VPWR VPWR _12789_/A sky130_fd_sc_hd__buf_1
XANTENNA_2 data_address[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14218_ _14506_/Q _14474_/Q _14442_/Q _14410_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14218_/X sky130_fd_sc_hd__mux4_2
XFILLER_99_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15198_ _08948_/X _15198_/D VGND VGND VPWR VPWR _15198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14149_ _14833_/Q _14865_/Q _14897_/Q _14929_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14149_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08710_ _08710_/A VGND VGND VPWR VPWR _08710_/X sky130_fd_sc_hd__clkbuf_2
X_09690_ _10827_/A VGND VGND VPWR VPWR _10431_/A sky130_fd_sc_hd__buf_1
XFILLER_27_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08641_ _15273_/Q _08637_/X _08511_/X _08638_/X VGND VGND VPWR VPWR _15273_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08572_ _08572_/A VGND VGND VPWR VPWR _08572_/X sky130_fd_sc_hd__clkbuf_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07454_ _07455_/A _13451_/X VGND VGND VPWR VPWR _15553_/D sky130_fd_sc_hd__and2_1
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07385_ _07491_/A _07385_/B VGND VGND VPWR VPWR _15594_/D sky130_fd_sc_hd__nor2_1
XFILLER_22_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09124_ _15147_/Q _09116_/X _08887_/X _09118_/X VGND VGND VPWR VPWR _15147_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09055_ _09055_/A VGND VGND VPWR VPWR _09117_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_136_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08006_ _08006_/A VGND VGND VPWR VPWR _08006_/X sky130_fd_sc_hd__buf_1
XFILLER_2_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09957_ _09972_/A VGND VGND VPWR VPWR _09957_/X sky130_fd_sc_hd__buf_1
XFILLER_58_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08908_ _08908_/A VGND VGND VPWR VPWR _08908_/X sky130_fd_sc_hd__clkbuf_1
X_09888_ _09888_/A VGND VGND VPWR VPWR _09908_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08839_ _09211_/A VGND VGND VPWR VPWR _08839_/X sky130_fd_sc_hd__buf_1
XFILLER_73_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11850_ _11850_/A VGND VGND VPWR VPWR _11907_/A sky130_fd_sc_hd__buf_1
XFILLER_122_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10801_ _14730_/Q _10797_/X _10799_/X _10800_/X VGND VGND VPWR VPWR _14730_/D sky130_fd_sc_hd__a22o_1
XFILLER_72_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11781_ _14472_/Q _11774_/X _11549_/X _11775_/X VGND VGND VPWR VPWR _14472_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13520_ _13519_/X _13060_/X _14336_/Q VGND VGND VPWR VPWR _13520_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10732_ _10764_/A VGND VGND VPWR VPWR _10732_/X sky130_fd_sc_hd__buf_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13451_ _13450_/X _13083_/X _14336_/Q VGND VGND VPWR VPWR _13451_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10663_ _10663_/A VGND VGND VPWR VPWR _10663_/X sky130_fd_sc_hd__buf_1
X_12402_ _15556_/Q VGND VGND VPWR VPWR _12415_/A sky130_fd_sc_hd__inv_2
X_13382_ _13384_/X _13383_/X _13415_/S VGND VGND VPWR VPWR _13382_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10594_ _14775_/Q _10584_/X _10349_/X _10585_/X VGND VGND VPWR VPWR _14775_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15121_ _09231_/X _15121_/D VGND VGND VPWR VPWR _15121_/Q sky130_fd_sc_hd__dfxtp_1
X_12333_ _12333_/A _12333_/B VGND VGND VPWR VPWR _12478_/A sky130_fd_sc_hd__or2_2
X_15052_ _09491_/X _15052_/D VGND VGND VPWR VPWR _15052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12264_ _12264_/A VGND VGND VPWR VPWR _12264_/X sky130_fd_sc_hd__buf_1
XFILLER_107_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14003_ _14687_/Q _15263_/Q _14751_/Q _14719_/Q _14055_/S0 _14057_/S1 VGND VGND VPWR
+ VPWR _14003_/X sky130_fd_sc_hd__mux4_2
X_11215_ _14624_/Q _11207_/X _11075_/X _11210_/X VGND VGND VPWR VPWR _14624_/D sky130_fd_sc_hd__a22o_1
X_12195_ _15569_/Q VGND VGND VPWR VPWR _12195_/X sky130_fd_sc_hd__clkbuf_2
X_11146_ _11151_/A VGND VGND VPWR VPWR _11146_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11077_ _11086_/A VGND VGND VPWR VPWR _11077_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10028_ _14925_/Q _10024_/X _10025_/X _10027_/X VGND VGND VPWR VPWR _14925_/D sky130_fd_sc_hd__a22o_1
X_14905_ _10105_/X _14905_/D VGND VGND VPWR VPWR _14905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14836_ _10362_/X _14836_/D VGND VGND VPWR VPWR _14836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14767_ _10621_/X _14767_/D VGND VGND VPWR VPWR _14767_/Q sky130_fd_sc_hd__dfxtp_1
X_11979_ _11981_/A VGND VGND VPWR VPWR _11979_/X sky130_fd_sc_hd__clkbuf_1
X_13718_ _14524_/Q _14492_/Q _14460_/Q _14428_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13718_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14698_ _10923_/X _14698_/D VGND VGND VPWR VPWR _14698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13649_ _13648_/X _07391_/Y _13649_/S VGND VGND VPWR VPWR _13649_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07170_ _07264_/B _07205_/A VGND VGND VPWR VPWR _07171_/B sky130_fd_sc_hd__or2_1
XFILLER_8_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15319_ _08417_/X _15319_/D VGND VGND VPWR VPWR _15319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09811_ _09823_/A VGND VGND VPWR VPWR _09812_/A sky130_fd_sc_hd__buf_1
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09742_ _14999_/Q _09736_/X _09589_/X _09737_/X VGND VGND VPWR VPWR _14999_/D sky130_fd_sc_hd__a22o_1
XFILLER_67_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09673_ _15016_/Q _09660_/X _09672_/X _09663_/X VGND VGND VPWR VPWR _15016_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08624_ _08635_/A VGND VGND VPWR VPWR _08633_/A sky130_fd_sc_hd__buf_1
XFILLER_82_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08555_ _08555_/A VGND VGND VPWR VPWR _08555_/X sky130_fd_sc_hd__buf_1
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07506_ _07506_/A _07506_/B VGND VGND VPWR VPWR _15518_/D sky130_fd_sc_hd__nor2_1
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08486_ _08486_/A VGND VGND VPWR VPWR _08524_/A sky130_fd_sc_hd__buf_1
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07437_ _07438_/A _13635_/X VGND VGND VPWR VPWR _15565_/D sky130_fd_sc_hd__and2_1
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07368_ _13154_/X _07363_/X _07506_/B _07354_/X _07367_/X VGND VGND VPWR VPWR _07370_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_109_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09107_ _09107_/A VGND VGND VPWR VPWR _09107_/X sky130_fd_sc_hd__buf_1
X_07299_ _14383_/Q VGND VGND VPWR VPWR _07505_/B sky130_fd_sc_hd__inv_2
X_09038_ _09038_/A VGND VGND VPWR VPWR _09038_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11000_ _11018_/A VGND VGND VPWR VPWR _11005_/A sky130_fd_sc_hd__buf_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12951_ _12951_/A _12951_/B _12951_/C VGND VGND VPWR VPWR _12951_/X sky130_fd_sc_hd__or3_4
XFILLER_46_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11902_ _14437_/Q _11895_/X _08091_/A _11896_/X VGND VGND VPWR VPWR _14437_/D sky130_fd_sc_hd__a22o_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15670_ _15672_/D _12986_/Y VGND VGND VPWR VPWR _15670_/Q sky130_fd_sc_hd__dlxtn_1
X_12882_ _13339_/X VGND VGND VPWR VPWR _12882_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_200 _13612_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_211 _13491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_222 _15491_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14621_ _11228_/X _14621_/D VGND VGND VPWR VPWR _14621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_233 _09886_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11833_ _11837_/A VGND VGND VPWR VPWR _11833_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_244 _11678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_255 _12753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14552_ _11478_/X _14552_/D VGND VGND VPWR VPWR _14552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11764_ _11783_/A VGND VGND VPWR VPWR _11764_/X sky130_fd_sc_hd__buf_1
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13503_ _13906_/X _13911_/X _13521_/S VGND VGND VPWR VPWR _13503_/X sky130_fd_sc_hd__mux2_1
X_10715_ _10721_/A VGND VGND VPWR VPWR _10715_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14483_ _11742_/X _14483_/D VGND VGND VPWR VPWR _14483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11695_ _11699_/A VGND VGND VPWR VPWR _11695_/X sky130_fd_sc_hd__clkbuf_1
X_13434_ _13676_/X _13681_/X _13521_/S VGND VGND VPWR VPWR _13434_/X sky130_fd_sc_hd__mux2_1
X_10646_ _10646_/A VGND VGND VPWR VPWR _10646_/X sky130_fd_sc_hd__buf_1
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13365_ _13367_/X _13366_/X _13415_/S VGND VGND VPWR VPWR _13365_/X sky130_fd_sc_hd__mux2_1
X_10577_ _14780_/Q _10575_/X _10328_/X _10576_/X VGND VGND VPWR VPWR _14780_/D sky130_fd_sc_hd__a22o_1
X_15104_ _09305_/X _15104_/D VGND VGND VPWR VPWR _15104_/Q sky130_fd_sc_hd__dfxtp_1
X_12316_ _12316_/A _12316_/B _12979_/B VGND VGND VPWR VPWR _12740_/A sky130_fd_sc_hd__or3_4
XFILLER_127_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13296_ _13297_/X _13315_/X _13415_/S VGND VGND VPWR VPWR _13296_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15035_ _09567_/X _15035_/D VGND VGND VPWR VPWR _15035_/Q sky130_fd_sc_hd__dfxtp_1
X_12247_ _12803_/A VGND VGND VPWR VPWR _12247_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12178_ _15540_/Q VGND VGND VPWR VPWR _12274_/A sky130_fd_sc_hd__inv_2
XFILLER_123_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11129_ _11137_/A VGND VGND VPWR VPWR _11129_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14819_ _10433_/X _14819_/D VGND VGND VPWR VPWR _14819_/Q sky130_fd_sc_hd__dfxtp_1
X_08340_ _14299_/Q _08340_/B _08778_/C VGND VGND VPWR VPWR _09521_/A sky130_fd_sc_hd__or3_1
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08271_ _08305_/A VGND VGND VPWR VPWR _08291_/A sky130_fd_sc_hd__clkbuf_2
X_07222_ _13102_/X _07220_/Y _07221_/X _07163_/B VGND VGND VPWR VPWR _15648_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07153_ _13094_/X VGND VGND VPWR VPWR _07286_/B sky130_fd_sc_hd__inv_2
XFILLER_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07986_ _07986_/A VGND VGND VPWR VPWR _07986_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09725_ _09731_/A VGND VGND VPWR VPWR _09725_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09656_ _10793_/A VGND VGND VPWR VPWR _10403_/A sky130_fd_sc_hd__buf_1
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08607_ _08617_/A VGND VGND VPWR VPWR _08607_/X sky130_fd_sc_hd__buf_1
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09587_ _09599_/A VGND VGND VPWR VPWR _09587_/X sky130_fd_sc_hd__clkbuf_1
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _14305_/Q VGND VGND VPWR VPWR _10827_/A sky130_fd_sc_hd__buf_1
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _08469_/A VGND VGND VPWR VPWR _08469_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10500_ _14802_/Q _10496_/X _10371_/X _10497_/X VGND VGND VPWR VPWR _14802_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11480_ _14552_/Q _11474_/X _11479_/X _11476_/X VGND VGND VPWR VPWR _14552_/D sky130_fd_sc_hd__a22o_1
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07523__1 _14313_/CLK VGND VGND VPWR VPWR _08294_/A sky130_fd_sc_hd__inv_2
XFILLER_109_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10431_ _10431_/A VGND VGND VPWR VPWR _10431_/X sky130_fd_sc_hd__buf_1
X_13150_ _12875_/B _12997_/Y _13152_/S VGND VGND VPWR VPWR _13150_/X sky130_fd_sc_hd__mux2_2
XFILLER_124_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10362_ _10370_/A VGND VGND VPWR VPWR _10362_/X sky130_fd_sc_hd__buf_1
XFILLER_124_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12101_ _15582_/Q VGND VGND VPWR VPWR _12101_/X sky130_fd_sc_hd__buf_1
X_13081_ _12609_/Y _15583_/Q _13090_/S VGND VGND VPWR VPWR _13081_/X sky130_fd_sc_hd__mux2_1
X_10293_ _10302_/A VGND VGND VPWR VPWR _10293_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12032_ _12024_/X _12029_/Y _13422_/X _12031_/X VGND VGND VPWR VPWR _12337_/A sky130_fd_sc_hd__o22a_2
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13983_ _14689_/Q _15265_/Q _14753_/Q _14721_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13983_/X sky130_fd_sc_hd__mux4_2
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12934_ _12958_/B _12930_/X _12805_/X _12812_/B _12933_/X VGND VGND VPWR VPWR _12934_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15653_ _15654_/CLK _15653_/D VGND VGND VPWR VPWR _15653_/Q sky130_fd_sc_hd__dfxtp_1
X_12865_ _12216_/Y _12864_/X _12216_/Y _12864_/X VGND VGND VPWR VPWR _12865_/Y sky130_fd_sc_hd__a2bb2oi_2
X_14604_ _11288_/X _14604_/D VGND VGND VPWR VPWR _14604_/Q sky130_fd_sc_hd__dfxtp_1
X_11816_ _11835_/A VGND VGND VPWR VPWR _11816_/X sky130_fd_sc_hd__buf_1
X_15584_ _15590_/CLK _15584_/D VGND VGND VPWR VPWR _15584_/Q sky130_fd_sc_hd__dfxtp_1
X_12796_ _12796_/A _13355_/X VGND VGND VPWR VPWR _12797_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14535_ _11551_/X _14535_/D VGND VGND VPWR VPWR _14535_/Q sky130_fd_sc_hd__dfxtp_1
X_11747_ _11751_/A VGND VGND VPWR VPWR _11747_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14466_ _11797_/X _14466_/D VGND VGND VPWR VPWR _14466_/Q sky130_fd_sc_hd__dfxtp_1
X_11678_ _11678_/A VGND VGND VPWR VPWR _11678_/X sky130_fd_sc_hd__clkbuf_1
X_13417_ _12838_/X _12847_/A _13418_/S VGND VGND VPWR VPWR _13417_/X sky130_fd_sc_hd__mux2_1
X_10629_ _10647_/A VGND VGND VPWR VPWR _10629_/X sky130_fd_sc_hd__buf_1
XFILLER_127_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14397_ _14397_/CLK instruction[22] VGND VGND VPWR VPWR _14397_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13348_ _13403_/X _13400_/X _13415_/S VGND VGND VPWR VPWR _13348_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13279_ _13278_/X _12345_/X _15565_/Q VGND VGND VPWR VPWR _13279_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15018_ _09659_/X _15018_/D VGND VGND VPWR VPWR _15018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07840_ _07786_/X _07678_/X _07849_/A _07703_/X _07681_/X VGND VGND VPWR VPWR _07846_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07771_ _07891_/A _07889_/B _07889_/A _07770_/X VGND VGND VPWR VPWR _07876_/A sky130_fd_sc_hd__a31o_1
XFILLER_37_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09510_ _09536_/A VGND VGND VPWR VPWR _09515_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09441_ _15067_/Q _09436_/X _09188_/X _09437_/X VGND VGND VPWR VPWR _15067_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09372_ _09372_/A VGND VGND VPWR VPWR _09381_/A sky130_fd_sc_hd__buf_1
X_08323_ _15336_/Q _08316_/X _08074_/X _08317_/X VGND VGND VPWR VPWR _15336_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08254_ _15356_/Q _08252_/X _07968_/X _08253_/X VGND VGND VPWR VPWR _15356_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07205_ _07205_/A VGND VGND VPWR VPWR _07205_/Y sky130_fd_sc_hd__inv_2
X_08185_ _08205_/A VGND VGND VPWR VPWR _08185_/X sky130_fd_sc_hd__buf_1
XFILLER_118_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07136_ _13108_/X VGND VGND VPWR VPWR _07267_/B sky130_fd_sc_hd__inv_2
XFILLER_118_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07969_ _07984_/A VGND VGND VPWR VPWR _07969_/X sky130_fd_sc_hd__buf_1
XFILLER_114_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09708_ _15009_/Q _09702_/X _09534_/X _09705_/X VGND VGND VPWR VPWR _15009_/D sky130_fd_sc_hd__a22o_1
X_10980_ _10984_/A VGND VGND VPWR VPWR _10980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09639_ _09647_/A VGND VGND VPWR VPWR _09639_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ _12578_/X _12642_/X _12644_/Y _12646_/X _12649_/X VGND VGND VPWR VPWR _12650_/Y
+ sky130_fd_sc_hd__o2111ai_4
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11601_ _11619_/A VGND VGND VPWR VPWR _11608_/A sky130_fd_sc_hd__buf_1
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ _12637_/A VGND VGND VPWR VPWR _12581_/X sky130_fd_sc_hd__buf_1
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14320_ _15599_/CLK _14320_/D VGND VGND VPWR VPWR _14320_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11532_ _11532_/A VGND VGND VPWR VPWR _11532_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ _14247_/X _14248_/X _14249_/X _14250_/X _14286_/S0 _14286_/S1 VGND VGND VPWR
+ VPWR _14251_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11463_ _11463_/A VGND VGND VPWR VPWR _11463_/X sky130_fd_sc_hd__buf_1
XFILLER_139_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13202_ _12590_/X _12577_/X _15561_/Q VGND VGND VPWR VPWR _13202_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10414_ _10422_/A VGND VGND VPWR VPWR _10414_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14182_ _15213_/Q _14541_/Q _14989_/Q _15405_/Q _14239_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14182_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11394_ _11414_/A VGND VGND VPWR VPWR _11394_/X sky130_fd_sc_hd__buf_1
XFILLER_151_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13133_ _12634_/X _13014_/Y _13152_/S VGND VGND VPWR VPWR _13133_/X sky130_fd_sc_hd__mux2_2
X_10345_ _14840_/Q _10339_/X _10344_/X _10341_/X VGND VGND VPWR VPWR _14840_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13064_ _12849_/Y _15566_/Q _13090_/S VGND VGND VPWR VPWR _13064_/X sky130_fd_sc_hd__mux2_1
X_10276_ _14857_/Q _10267_/X _10042_/X _10268_/X VGND VGND VPWR VPWR _14857_/D sky130_fd_sc_hd__a22o_1
X_12015_ _12017_/A VGND VGND VPWR VPWR _12015_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13966_ _13962_/X _13963_/X _13964_/X _13965_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13966_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12917_ _12791_/X _12195_/X _12775_/A _12788_/X VGND VGND VPWR VPWR _12919_/C sky130_fd_sc_hd__o22a_1
XFILLER_74_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13897_ _14634_/Q _14602_/Q _14570_/Q _15370_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13897_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15636_ _15668_/CLK _15636_/D VGND VGND VPWR VPWR pc[31] sky130_fd_sc_hd__dfxtp_4
X_12848_ _13309_/X _12782_/X _12821_/A _12846_/X _12847_/X VGND VGND VPWR VPWR _12848_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15567_ _15578_/CLK _15567_/D VGND VGND VPWR VPWR _15567_/Q sky130_fd_sc_hd__dfxtp_1
X_12779_ _12779_/A VGND VGND VPWR VPWR _12785_/B sky130_fd_sc_hd__buf_1
XFILLER_42_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14518_ _11620_/X _14518_/D VGND VGND VPWR VPWR _14518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15498_ _15498_/CLK _15498_/D VGND VGND VPWR VPWR wdata[24] sky130_fd_sc_hd__dfxtp_4
XFILLER_147_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14449_ _11862_/X _14449_/D VGND VGND VPWR VPWR _14449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09990_ _09990_/A VGND VGND VPWR VPWR _09990_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08941_ _08941_/A VGND VGND VPWR VPWR _09005_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08872_ _08882_/A VGND VGND VPWR VPWR _08872_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07823_ _07786_/X _07686_/X _07778_/C _07832_/B _07695_/A VGND VGND VPWR VPWR _07830_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07754_ _07754_/A _15596_/Q VGND VGND VPWR VPWR _07754_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07685_ _07653_/A _07678_/X _07681_/X _07684_/X VGND VGND VPWR VPWR _07779_/A sky130_fd_sc_hd__o211a_1
XFILLER_92_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09424_ _09485_/A VGND VGND VPWR VPWR _09445_/A sky130_fd_sc_hd__clkbuf_2
X_09355_ _09361_/A VGND VGND VPWR VPWR _09355_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08306_ _08325_/A VGND VGND VPWR VPWR _08306_/X sky130_fd_sc_hd__buf_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09286_ _09289_/A VGND VGND VPWR VPWR _09286_/X sky130_fd_sc_hd__clkbuf_1
X_08237_ _15360_/Q _08227_/X _07944_/X _08230_/X VGND VGND VPWR VPWR _15360_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08168_ _15378_/Q _08164_/X _08021_/X _08165_/X VGND VGND VPWR VPWR _15378_/D sky130_fd_sc_hd__a22o_1
XFILLER_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07119_ _15512_/Q VGND VGND VPWR VPWR _12030_/C sky130_fd_sc_hd__inv_2
XFILLER_107_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08099_ _08099_/A VGND VGND VPWR VPWR _08099_/X sky130_fd_sc_hd__clkbuf_2
X_10130_ _10132_/A VGND VGND VPWR VPWR _10130_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10061_ _10064_/A VGND VGND VPWR VPWR _10061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13820_ _14962_/Q _15058_/Q _15026_/Q _15090_/Q _13860_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13820_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13751_ _13747_/X _13748_/X _13749_/X _13750_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13751_/X sky130_fd_sc_hd__mux4_1
X_10963_ _11024_/A VGND VGND VPWR VPWR _10985_/A sky130_fd_sc_hd__clkbuf_2
X_12702_ _12784_/A VGND VGND VPWR VPWR _12758_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_44_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13682_ _15231_/Q _14559_/Q _15007_/Q _15423_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13682_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10894_ _10904_/A VGND VGND VPWR VPWR _10894_/X sky130_fd_sc_hd__buf_1
X_15421_ _07961_/X _15421_/D VGND VGND VPWR VPWR _15421_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12633_ _12428_/X _12612_/Y _12625_/X _12629_/X _12632_/Y VGND VGND VPWR VPWR _12633_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_34_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15352_ _08266_/X _15352_/D VGND VGND VPWR VPWR _15352_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12564_ _14391_/Q _14390_/Q _14389_/Q _14388_/Q VGND VGND VPWR VPWR _12565_/C sky130_fd_sc_hd__or4_4
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ _15469_/CLK _15470_/Q VGND VGND VPWR VPWR _14303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11515_ _11515_/A VGND VGND VPWR VPWR _11515_/X sky130_fd_sc_hd__buf_1
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15283_ _08606_/X _15283_/D VGND VGND VPWR VPWR _15283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12495_ _12495_/A VGND VGND VPWR VPWR _12951_/A sky130_fd_sc_hd__buf_1
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14234_ _15176_/Q _15144_/Q _14760_/Q _14792_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14234_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11446_ _11446_/A VGND VGND VPWR VPWR _11526_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14165_ _15119_/Q _15343_/Q _15311_/Q _15279_/Q _14238_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14165_/X sky130_fd_sc_hd__mux4_2
X_11377_ _11407_/A VGND VGND VPWR VPWR _11398_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13116_ _15662_/Q data_address[27] _15667_/Q VGND VGND VPWR VPWR _13116_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10328_ _10328_/A VGND VGND VPWR VPWR _10328_/X sky130_fd_sc_hd__buf_1
X_14096_ _14092_/X _14093_/X _14094_/X _14095_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14096_/X sky130_fd_sc_hd__mux4_2
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13047_ wdata[20] rdata[20] _13057_/S VGND VGND VPWR VPWR _14324_/D sky130_fd_sc_hd__mux2_1
X_10259_ _10281_/A VGND VGND VPWR VPWR _10259_/X sky130_fd_sc_hd__buf_1
XFILLER_94_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14998_ _09744_/X _14998_/D VGND VGND VPWR VPWR _14998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13949_ _14821_/Q _14853_/Q _14885_/Q _14917_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13949_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07470_ _07472_/A _13484_/X VGND VGND VPWR VPWR _15542_/D sky130_fd_sc_hd__and2_1
XFILLER_61_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15619_ _15621_/CLK _15619_/D VGND VGND VPWR VPWR pc[14] sky130_fd_sc_hd__dfxtp_2
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09140_ _09144_/A VGND VGND VPWR VPWR _09140_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09071_ _15163_/Q _09065_/X _08817_/X _09066_/X VGND VGND VPWR VPWR _15163_/D sky130_fd_sc_hd__a22o_1
X_08022_ _15410_/Q _08014_/X _08021_/X _08017_/X VGND VGND VPWR VPWR _15410_/D sky130_fd_sc_hd__a22o_1
XFILLER_135_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09973_ _10340_/A VGND VGND VPWR VPWR _09973_/X sky130_fd_sc_hd__buf_1
X_08924_ _11062_/B VGND VGND VPWR VPWR _10294_/A sky130_fd_sc_hd__buf_1
XFILLER_69_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08855_ _08855_/A VGND VGND VPWR VPWR _08855_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07806_ _07659_/X _07671_/X _07805_/Y VGND VGND VPWR VPWR _07807_/A sky130_fd_sc_hd__o21ai_1
X_08786_ _08786_/A VGND VGND VPWR VPWR _08786_/X sky130_fd_sc_hd__buf_1
XFILLER_44_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07737_ _07874_/A _07875_/A VGND VGND VPWR VPWR _07772_/C sky130_fd_sc_hd__nand2_1
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07668_ _07668_/A VGND VGND VPWR VPWR _07668_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09407_ _09407_/A VGND VGND VPWR VPWR _09407_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07599_ _07599_/A _13068_/X VGND VGND VPWR VPWR _15483_/D sky130_fd_sc_hd__and2_1
XFILLER_41_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09338_ _09340_/A VGND VGND VPWR VPWR _09338_/X sky130_fd_sc_hd__clkbuf_1
X_09269_ _09269_/A VGND VGND VPWR VPWR _09278_/A sky130_fd_sc_hd__buf_1
X_11300_ _14600_/Q _11294_/X _11183_/X _11295_/X VGND VGND VPWR VPWR _14600_/D sky130_fd_sc_hd__a22o_1
X_12280_ _12692_/A VGND VGND VPWR VPWR _12693_/A sky130_fd_sc_hd__inv_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11231_ _11237_/A VGND VGND VPWR VPWR _11231_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11162_ _11162_/A VGND VGND VPWR VPWR _11188_/A sky130_fd_sc_hd__buf_1
XFILLER_96_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10113_ _10143_/A VGND VGND VPWR VPWR _10134_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11093_ _11098_/A VGND VGND VPWR VPWR _11093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10044_ _10044_/A VGND VGND VPWR VPWR _10067_/A sky130_fd_sc_hd__clkbuf_2
X_14921_ _10041_/X _14921_/D VGND VGND VPWR VPWR _14921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14852_ _10288_/X _14852_/D VGND VGND VPWR VPWR _14852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13803_ _14675_/Q _15251_/Q _14739_/Q _14707_/Q _13918_/S0 _13860_/S1 VGND VGND VPWR
+ VPWR _13803_/X sky130_fd_sc_hd__mux4_2
X_14783_ _10561_/X _14783_/D VGND VGND VPWR VPWR _14783_/Q sky130_fd_sc_hd__dfxtp_1
X_11995_ _12001_/A VGND VGND VPWR VPWR _11995_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13734_ _15194_/Q _15162_/Q _14778_/Q _14810_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13734_/X sky130_fd_sc_hd__mux4_2
X_10946_ _10948_/A VGND VGND VPWR VPWR _10946_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13665_ _15137_/Q _15361_/Q _15329_/Q _15297_/Q _13740_/S0 _07541_/A VGND VGND VPWR
+ VPWR _13665_/X sky130_fd_sc_hd__mux4_1
X_10877_ _10879_/A VGND VGND VPWR VPWR _10877_/X sky130_fd_sc_hd__clkbuf_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12616_ _12616_/A VGND VGND VPWR VPWR _12616_/X sky130_fd_sc_hd__clkbuf_2
X_15404_ _08052_/X _15404_/D VGND VGND VPWR VPWR _15404_/Q sky130_fd_sc_hd__dfxtp_1
X_13596_ _14156_/X _14161_/X _13648_/S VGND VGND VPWR VPWR _13596_/X sky130_fd_sc_hd__mux2_2
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15335_ _08324_/X _15335_/D VGND VGND VPWR VPWR _15335_/Q sky130_fd_sc_hd__dfxtp_1
X_12547_ data_address[1] VGND VGND VPWR VPWR _12556_/A sky130_fd_sc_hd__buf_1
XFILLER_129_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15266_ _08659_/X _15266_/D VGND VGND VPWR VPWR _15266_/Q sky130_fd_sc_hd__dfxtp_1
X_12478_ _12478_/A VGND VGND VPWR VPWR _12784_/A sky130_fd_sc_hd__buf_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_3 data_address[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14217_ _14634_/Q _14602_/Q _14570_/Q _15370_/Q _14268_/S0 _07379_/A VGND VGND VPWR
+ VPWR _14217_/X sky130_fd_sc_hd__mux4_1
X_11429_ _11446_/A VGND VGND VPWR VPWR _11430_/A sky130_fd_sc_hd__buf_1
X_15197_ _08950_/X _15197_/D VGND VGND VPWR VPWR _15197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14148_ _14513_/Q _14481_/Q _14449_/Q _14417_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14148_/X sky130_fd_sc_hd__mux4_2
XFILLER_125_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14079_ _14840_/Q _14872_/Q _14904_/Q _14936_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14079_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08640_ _08642_/A VGND VGND VPWR VPWR _08640_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08571_ _15294_/Q _08565_/X _08377_/X _08568_/X VGND VGND VPWR VPWR _15294_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_46_clk _14315_/CLK VGND VGND VPWR VPWR _15601_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07522_ _07641_/A _14371_/Q VGND VGND VPWR VPWR _15507_/D sky130_fd_sc_hd__or2_1
X_07453_ _07455_/A _13448_/X VGND VGND VPWR VPWR _15554_/D sky130_fd_sc_hd__and2_1
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07384_ _07496_/A VGND VGND VPWR VPWR _07491_/A sky130_fd_sc_hd__buf_1
X_09123_ _09125_/A VGND VGND VPWR VPWR _09123_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09054_ _09075_/A VGND VGND VPWR VPWR _09054_/X sky130_fd_sc_hd__buf_1
X_08005_ _14322_/Q VGND VGND VPWR VPWR _08006_/A sky130_fd_sc_hd__buf_1
XFILLER_144_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09956_ _09961_/A VGND VGND VPWR VPWR _09956_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08907_ _15207_/Q _08904_/X _08905_/X _08906_/X VGND VGND VPWR VPWR _15207_/D sky130_fd_sc_hd__a22o_1
X_09887_ _09907_/A VGND VGND VPWR VPWR _09887_/X sky130_fd_sc_hd__buf_1
XFILLER_73_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08838_ _08864_/A VGND VGND VPWR VPWR _08838_/X sky130_fd_sc_hd__buf_1
XFILLER_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08769_ _15237_/Q _08762_/X _08535_/X _08763_/X VGND VGND VPWR VPWR _15237_/D sky130_fd_sc_hd__a22o_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_37_clk _14397_/CLK VGND VGND VPWR VPWR _15578_/CLK sky130_fd_sc_hd__clkbuf_16
X_10800_ _10815_/A VGND VGND VPWR VPWR _10800_/X sky130_fd_sc_hd__buf_1
X_11780_ _11782_/A VGND VGND VPWR VPWR _11780_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10731_ _10779_/A VGND VGND VPWR VPWR _10764_/A sky130_fd_sc_hd__buf_1
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13450_ _13449_/X rdata[24] _13516_/S VGND VGND VPWR VPWR _13450_/X sky130_fd_sc_hd__mux2_2
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10662_ _10680_/A VGND VGND VPWR VPWR _10663_/A sky130_fd_sc_hd__buf_1
XFILLER_139_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12401_ _12401_/A VGND VGND VPWR VPWR _12410_/A sky130_fd_sc_hd__buf_1
X_13381_ _12785_/A _12762_/X _13418_/S VGND VGND VPWR VPWR _13381_/X sky130_fd_sc_hd__mux2_1
X_10593_ _10595_/A VGND VGND VPWR VPWR _10593_/X sky130_fd_sc_hd__clkbuf_1
X_15120_ _09234_/X _15120_/D VGND VGND VPWR VPWR _15120_/Q sky130_fd_sc_hd__dfxtp_1
X_12332_ _12319_/X _12323_/X _12328_/X _12904_/A VGND VGND VPWR VPWR _12342_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15051_ _09493_/X _15051_/D VGND VGND VPWR VPWR _15051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12263_ _12264_/A _12265_/A _12798_/A _12799_/A VGND VGND VPWR VPWR _12263_/X sky130_fd_sc_hd__and4_1
XFILLER_142_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14002_ _15231_/Q _14559_/Q _15007_/Q _15423_/Q _14395_/Q _14057_/S1 VGND VGND VPWR
+ VPWR _14002_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11214_ _11214_/A VGND VGND VPWR VPWR _11214_/X sky130_fd_sc_hd__clkbuf_1
X_12194_ _15537_/Q VGND VGND VPWR VPWR _12774_/A sky130_fd_sc_hd__inv_2
XFILLER_150_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11145_ _14641_/Q _11133_/X _11144_/X _11135_/X VGND VGND VPWR VPWR _14641_/D sky130_fd_sc_hd__a22o_1
XFILLER_122_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11076_ _14656_/Q _11064_/X _11075_/X _11068_/X VGND VGND VPWR VPWR _14656_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10027_ _10052_/A VGND VGND VPWR VPWR _10027_/X sky130_fd_sc_hd__buf_1
X_14904_ _10109_/X _14904_/D VGND VGND VPWR VPWR _14904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14835_ _10365_/X _14835_/D VGND VGND VPWR VPWR _14835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_clk _14397_/CLK VGND VGND VPWR VPWR _15621_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11978_ _14416_/Q _11976_/X _08031_/A _11977_/X VGND VGND VPWR VPWR _14416_/D sky130_fd_sc_hd__a22o_1
X_14766_ _10623_/X _14766_/D VGND VGND VPWR VPWR _14766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10929_ _10929_/A VGND VGND VPWR VPWR _10929_/X sky130_fd_sc_hd__clkbuf_1
X_13717_ _14652_/Q _14620_/Q _14588_/Q _15388_/Q _13737_/S0 _13740_/S1 VGND VGND VPWR
+ VPWR _13717_/X sky130_fd_sc_hd__mux4_2
X_14697_ _10927_/X _14697_/D VGND VGND VPWR VPWR _14697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13648_ _14286_/X _14291_/X _13648_/S VGND VGND VPWR VPWR _13648_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13579_ _13578_/X _13077_/X _14337_/Q VGND VGND VPWR VPWR _13579_/X sky130_fd_sc_hd__mux2_1
X_15318_ _08422_/X _15318_/D VGND VGND VPWR VPWR _15318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15249_ _08729_/X _15249_/D VGND VGND VPWR VPWR _15249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09810_ _10294_/A _09810_/B VGND VGND VPWR VPWR _09823_/A sky130_fd_sc_hd__or2_2
XFILLER_98_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09741_ _09741_/A VGND VGND VPWR VPWR _09741_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09672_ _10415_/A VGND VGND VPWR VPWR _09672_/X sky130_fd_sc_hd__buf_1
XFILLER_39_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08623_ _15278_/Q _08617_/X _08478_/X _08618_/X VGND VGND VPWR VPWR _15278_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clk _14397_/CLK VGND VGND VPWR VPWR _15566_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08554_ _08566_/A VGND VGND VPWR VPWR _08555_/A sky130_fd_sc_hd__buf_1
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07505_ _07506_/A _07505_/B VGND VGND VPWR VPWR _15519_/D sky130_fd_sc_hd__nor2_1
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08485_ _09250_/A VGND VGND VPWR VPWR _08485_/X sky130_fd_sc_hd__buf_1
XFILLER_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07436_ _07438_/A _13631_/X VGND VGND VPWR VPWR _15566_/D sky130_fd_sc_hd__and2_1
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07367_ _07508_/B _07356_/X _12573_/A _07308_/X VGND VGND VPWR VPWR _07367_/X sky130_fd_sc_hd__o22a_1
X_09106_ _09106_/A VGND VGND VPWR VPWR _09106_/X sky130_fd_sc_hd__buf_1
XFILLER_136_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07298_ _07363_/A VGND VGND VPWR VPWR _07298_/X sky130_fd_sc_hd__clkbuf_2
X_09037_ _15171_/Q _08929_/A _08919_/X _08932_/A VGND VGND VPWR VPWR _15171_/D sky130_fd_sc_hd__a22o_1
XFILLER_144_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09939_ _14944_/Q _09927_/X _09938_/X _09931_/X VGND VGND VPWR VPWR _14944_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12950_ _12588_/X _12591_/X _12959_/D _12942_/X _12949_/X VGND VGND VPWR VPWR _12950_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_18_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11901_ _11905_/A VGND VGND VPWR VPWR _11901_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12881_ _12874_/Y _12876_/X _12663_/X _12877_/X _12880_/X VGND VGND VPWR VPWR _12881_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_45_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_201 _13590_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_212 _13492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_223 _15506_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11832_ _14458_/Q _11825_/X _07978_/A _11826_/X VGND VGND VPWR VPWR _14458_/D sky130_fd_sc_hd__a22o_1
X_14620_ _11231_/X _14620_/D VGND VGND VPWR VPWR _14620_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_234 _09846_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_245 _11907_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_256 _12753_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14551_ _11483_/X _14551_/D VGND VGND VPWR VPWR _14551_/Q sky130_fd_sc_hd__dfxtp_1
X_11763_ _11763_/A VGND VGND VPWR VPWR _11783_/A sky130_fd_sc_hd__buf_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10714_ _14746_/Q _10701_/X _10713_/X _10704_/X VGND VGND VPWR VPWR _14746_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13502_ _13501_/X _13066_/X _14336_/Q VGND VGND VPWR VPWR _13502_/X sky130_fd_sc_hd__mux2_1
X_14482_ _11747_/X _14482_/D VGND VGND VPWR VPWR _14482_/Q sky130_fd_sc_hd__dfxtp_1
X_11694_ _11716_/A VGND VGND VPWR VPWR _11699_/A sky130_fd_sc_hd__buf_1
X_13433_ _13432_/X _13089_/X _14336_/Q VGND VGND VPWR VPWR _13433_/X sky130_fd_sc_hd__mux2_1
X_10645_ _10645_/A VGND VGND VPWR VPWR _10645_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13364_ _12480_/B _12492_/X _13418_/S VGND VGND VPWR VPWR _13364_/X sky130_fd_sc_hd__mux2_1
X_10576_ _10585_/A VGND VGND VPWR VPWR _10576_/X sky130_fd_sc_hd__buf_1
XFILLER_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12315_ _12315_/A VGND VGND VPWR VPWR _12699_/A sky130_fd_sc_hd__buf_1
X_15103_ _09308_/X _15103_/D VGND VGND VPWR VPWR _15103_/Q sky130_fd_sc_hd__dfxtp_1
X_13295_ _12835_/Y _13338_/X _13408_/S VGND VGND VPWR VPWR _13295_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15034_ _09572_/X _15034_/D VGND VGND VPWR VPWR _15034_/Q sky130_fd_sc_hd__dfxtp_1
X_12246_ _12246_/A _12246_/B VGND VGND VPWR VPWR _12803_/A sky130_fd_sc_hd__or2_1
XFILLER_108_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12177_ _12162_/Y _12685_/A _12684_/A VGND VGND VPWR VPWR _12177_/Y sky130_fd_sc_hd__nand3b_2
X_11128_ _11128_/A VGND VGND VPWR VPWR _11137_/A sky130_fd_sc_hd__buf_2
X_11059_ _14659_/Q _10951_/A _10832_/X _10954_/A VGND VGND VPWR VPWR _14659_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14818_ _10437_/X _14818_/D VGND VGND VPWR VPWR _14818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14749_ _10696_/X _14749_/D VGND VGND VPWR VPWR _14749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08270_ _08270_/A VGND VGND VPWR VPWR _08270_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07221_ _07221_/A VGND VGND VPWR VPWR _07221_/X sky130_fd_sc_hd__buf_1
XFILLER_146_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07152_ _13093_/X VGND VGND VPWR VPWR _07242_/A sky130_fd_sc_hd__inv_2
XFILLER_146_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clkbuf_opt_8_clk/A VGND VGND VPWR VPWR _14313_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07985_ _15417_/Q _07981_/X _07983_/X _07984_/X VGND VGND VPWR VPWR _15417_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09724_ _09724_/A VGND VGND VPWR VPWR _09731_/A sky130_fd_sc_hd__buf_1
XFILLER_28_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09655_ _09665_/A VGND VGND VPWR VPWR _09655_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08606_ _08612_/A VGND VGND VPWR VPWR _08606_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09586_ _09586_/A VGND VGND VPWR VPWR _09599_/A sky130_fd_sc_hd__buf_2
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08537_ _08542_/A VGND VGND VPWR VPWR _08537_/X sky130_fd_sc_hd__clkbuf_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ _15312_/Q _08463_/X _08466_/X _08467_/X VGND VGND VPWR VPWR _15312_/D sky130_fd_sc_hd__a22o_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07419_ _07419_/A _13591_/X VGND VGND VPWR VPWR _15576_/D sky130_fd_sc_hd__and2_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08399_ _08411_/A VGND VGND VPWR VPWR _08399_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_10430_ _10433_/A VGND VGND VPWR VPWR _10430_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07523__2 _14313_/CLK VGND VGND VPWR VPWR _07524_/A sky130_fd_sc_hd__inv_2
XFILLER_148_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10361_ _10373_/A VGND VGND VPWR VPWR _10370_/A sky130_fd_sc_hd__buf_1
XFILLER_152_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12100_ _12109_/A VGND VGND VPWR VPWR _12610_/A sky130_fd_sc_hd__buf_1
XFILLER_124_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13080_ _12624_/Y _15582_/Q _13090_/S VGND VGND VPWR VPWR _13080_/X sky130_fd_sc_hd__mux2_1
X_10292_ _14851_/Q _10183_/A _10065_/X _10186_/A VGND VGND VPWR VPWR _14851_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12031_ _12031_/A VGND VGND VPWR VPWR _12031_/X sky130_fd_sc_hd__buf_1
XFILLER_3_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13982_ _15233_/Q _14561_/Q _15009_/Q _15425_/Q _14060_/S0 _14060_/S1 VGND VGND VPWR
+ VPWR _13982_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12933_ _12933_/A _12933_/B VGND VGND VPWR VPWR _12933_/X sky130_fd_sc_hd__or2_1
XFILLER_58_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15652_ _15652_/CLK _15652_/D VGND VGND VPWR VPWR _15652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12864_ _12875_/B _12220_/A _12228_/A _12863_/Y VGND VGND VPWR VPWR _12864_/X sky130_fd_sc_hd__o22a_1
X_14603_ _11290_/X _14603_/D VGND VGND VPWR VPWR _14603_/Q sky130_fd_sc_hd__dfxtp_1
X_11815_ _11876_/A VGND VGND VPWR VPWR _11835_/A sky130_fd_sc_hd__buf_2
X_12795_ _13280_/X _12707_/X _12790_/X _12793_/Y _12794_/X VGND VGND VPWR VPWR _12795_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_15583_ _15591_/CLK _15583_/D VGND VGND VPWR VPWR _15583_/Q sky130_fd_sc_hd__dfxtp_1
X_11746_ _11746_/A VGND VGND VPWR VPWR _11751_/A sky130_fd_sc_hd__buf_1
X_14534_ _11556_/X _14534_/D VGND VGND VPWR VPWR _14534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14465_ _11805_/X _14465_/D VGND VGND VPWR VPWR _14465_/Q sky130_fd_sc_hd__dfxtp_1
X_11677_ _14502_/Q _11673_/X _11557_/X _11674_/X VGND VGND VPWR VPWR _14502_/D sky130_fd_sc_hd__a22o_1
XFILLER_146_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13416_ _12820_/X _12812_/A _13418_/S VGND VGND VPWR VPWR _13416_/X sky130_fd_sc_hd__mux2_1
X_10628_ _10628_/A VGND VGND VPWR VPWR _10647_/A sky130_fd_sc_hd__clkbuf_2
X_14396_ _15666_/CLK instruction[21] VGND VGND VPWR VPWR _14396_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13347_ _13349_/X _13348_/X _13408_/S VGND VGND VPWR VPWR _13347_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10559_ _10561_/A VGND VGND VPWR VPWR _10559_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13278_ _13375_/X _13368_/X _13393_/S VGND VGND VPWR VPWR _13278_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12229_ _15531_/Q VGND VGND VPWR VPWR _12929_/B sky130_fd_sc_hd__buf_1
X_15017_ _09665_/X _15017_/D VGND VGND VPWR VPWR _15017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07770_ _07743_/Y _15599_/Q _07769_/X _07739_/X _07740_/X VGND VGND VPWR VPWR _07770_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09440_ _09444_/A VGND VGND VPWR VPWR _09440_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09371_ _15086_/Q _09365_/X _09245_/X _09366_/X VGND VGND VPWR VPWR _15086_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08322_ _08324_/A VGND VGND VPWR VPWR _08322_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08253_ _08262_/A VGND VGND VPWR VPWR _08253_/X sky130_fd_sc_hd__buf_1
XFILLER_119_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07204_ _07263_/B _07171_/B _07200_/X _07202_/Y VGND VGND VPWR VPWR _15657_/D sky130_fd_sc_hd__a211oi_2
XFILLER_137_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08184_ _08184_/A VGND VGND VPWR VPWR _08205_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07135_ _13109_/X VGND VGND VPWR VPWR _07265_/B sky130_fd_sc_hd__inv_2
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07968_ _07968_/A VGND VGND VPWR VPWR _07968_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09707_ _09709_/A VGND VGND VPWR VPWR _09707_/X sky130_fd_sc_hd__clkbuf_1
X_07899_ _07765_/Y _07752_/Y _07893_/X _07895_/X VGND VGND VPWR VPWR _15431_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09638_ _15022_/Q _09625_/X _09637_/X _09628_/X VGND VGND VPWR VPWR _15022_/D sky130_fd_sc_hd__a22o_1
XFILLER_43_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09569_ _10332_/A VGND VGND VPWR VPWR _09569_/X sky130_fd_sc_hd__buf_1
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _11630_/A VGND VGND VPWR VPWR _11619_/A sky130_fd_sc_hd__clkbuf_4
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _12580_/A VGND VGND VPWR VPWR _12625_/A sky130_fd_sc_hd__buf_1
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ _14541_/Q _11527_/X _11528_/X _11530_/X VGND VGND VPWR VPWR _14541_/D sky130_fd_sc_hd__a22o_1
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _14951_/Q _15047_/Q _15015_/Q _15079_/Q _07387_/A _07379_/A VGND VGND VPWR
+ VPWR _14250_/X sky130_fd_sc_hd__mux4_2
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11462_ _11474_/A VGND VGND VPWR VPWR _11462_/X sky130_fd_sc_hd__buf_1
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ _13202_/X _13212_/X _15562_/Q VGND VGND VPWR VPWR _13201_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10413_ _10413_/A VGND VGND VPWR VPWR _10422_/A sky130_fd_sc_hd__buf_1
X_14181_ _14177_/X _14178_/X _14179_/X _14180_/X _14397_/Q _14266_/S1 VGND VGND VPWR
+ VPWR _14181_/X sky130_fd_sc_hd__mux4_1
X_11393_ _11393_/A VGND VGND VPWR VPWR _11414_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13132_ _12611_/X _13015_/Y _13152_/S VGND VGND VPWR VPWR _13132_/X sky130_fd_sc_hd__mux2_2
X_10344_ _10344_/A VGND VGND VPWR VPWR _10344_/X sky130_fd_sc_hd__buf_1
XFILLER_152_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13063_ _12858_/Y _15565_/Q _13090_/S VGND VGND VPWR VPWR _13063_/X sky130_fd_sc_hd__mux2_2
X_10275_ _10279_/A VGND VGND VPWR VPWR _10275_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12014_ _14404_/Q _11912_/A _08095_/A _11915_/A VGND VGND VPWR VPWR _14404_/D sky130_fd_sc_hd__a22o_1
XFILLER_105_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13965_ _15107_/Q _15331_/Q _15299_/Q _15267_/Q _07542_/A _07541_/A VGND VGND VPWR
+ VPWR _13965_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12916_ _12752_/X _12179_/X _12754_/A _12755_/A VGND VGND VPWR VPWR _12937_/A sky130_fd_sc_hd__o22a_1
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13896_ _13892_/X _13893_/X _13894_/X _13895_/X _14401_/Q _13946_/S1 VGND VGND VPWR
+ VPWR _13896_/X sky130_fd_sc_hd__mux4_2
XFILLER_34_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15635_ _15654_/CLK _15635_/D VGND VGND VPWR VPWR pc[30] sky130_fd_sc_hd__dfxtp_4
X_12847_ _12847_/A _12847_/B _12847_/C VGND VGND VPWR VPWR _12847_/X sky130_fd_sc_hd__or3_1
XFILLER_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15566_ _15566_/CLK _15566_/D VGND VGND VPWR VPWR _15566_/Q sky130_fd_sc_hd__dfxtp_1
X_12778_ _15538_/Q VGND VGND VPWR VPWR _12778_/X sky130_fd_sc_hd__buf_1
XFILLER_15_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14517_ _11626_/X _14517_/D VGND VGND VPWR VPWR _14517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11729_ _11731_/A VGND VGND VPWR VPWR _11729_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15497_ _15590_/CLK _15497_/D VGND VGND VPWR VPWR wdata[23] sky130_fd_sc_hd__dfxtp_2
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14448_ _11864_/X _14448_/D VGND VGND VPWR VPWR _14448_/Q sky130_fd_sc_hd__dfxtp_1
X_14379_ _14379_/CLK instruction[8] VGND VGND VPWR VPWR _14379_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08940_ _08950_/A VGND VGND VPWR VPWR _08940_/X sky130_fd_sc_hd__clkbuf_1
X_08871_ _08885_/A VGND VGND VPWR VPWR _08882_/A sky130_fd_sc_hd__buf_2
XFILLER_111_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07822_ _07822_/A VGND VGND VPWR VPWR _07832_/B sky130_fd_sc_hd__inv_2
XFILLER_97_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07753_ _13149_/X VGND VGND VPWR VPWR _07754_/A sky130_fd_sc_hd__inv_2
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07684_ _07682_/X _07683_/X _07682_/X _13133_/X VGND VGND VPWR VPWR _07684_/X sky130_fd_sc_hd__o22a_1
XFILLER_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09423_ _09423_/A VGND VGND VPWR VPWR _09485_/A sky130_fd_sc_hd__buf_2
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09354_ _09372_/A VGND VGND VPWR VPWR _09361_/A sky130_fd_sc_hd__buf_1
XFILLER_52_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08305_ _08305_/A VGND VGND VPWR VPWR _08325_/A sky130_fd_sc_hd__buf_1
X_09285_ _15109_/Q _09274_/X _09284_/X _09276_/X VGND VGND VPWR VPWR _15109_/D sky130_fd_sc_hd__a22o_1
XFILLER_138_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08236_ _08238_/A VGND VGND VPWR VPWR _08236_/X sky130_fd_sc_hd__clkbuf_1
X_08167_ _08169_/A VGND VGND VPWR VPWR _08167_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_07118_ _12040_/A VGND VGND VPWR VPWR _07634_/B sky130_fd_sc_hd__inv_2
XFILLER_134_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08098_ _14304_/Q VGND VGND VPWR VPWR _08099_/A sky130_fd_sc_hd__buf_1
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10060_ _14917_/Q _10050_/X _10059_/X _10052_/X VGND VGND VPWR VPWR _14917_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10962_ _10962_/A VGND VGND VPWR VPWR _11024_/A sky130_fd_sc_hd__buf_4
X_13750_ _14969_/Q _15065_/Q _15033_/Q _15097_/Q _13963_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13750_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12701_ _12706_/A VGND VGND VPWR VPWR _12701_/X sky130_fd_sc_hd__buf_1
XFILLER_44_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10893_ _10899_/A VGND VGND VPWR VPWR _10893_/X sky130_fd_sc_hd__clkbuf_1
X_13681_ _13677_/X _13678_/X _13679_/X _13680_/X _07533_/A _14402_/Q VGND VGND VPWR
+ VPWR _13681_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15420_ _07965_/X _15420_/D VGND VGND VPWR VPWR _15420_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12632_ _12632_/A _12632_/B VGND VGND VPWR VPWR _12632_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _12563_/A _14383_/Q _12563_/C VGND VGND VPWR VPWR _13157_/S sky130_fd_sc_hd__and3_2
X_15351_ _08268_/X _15351_/D VGND VGND VPWR VPWR _15351_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11514_ _11514_/A VGND VGND VPWR VPWR _11514_/X sky130_fd_sc_hd__buf_1
X_14302_ _15469_/CLK _15469_/Q VGND VGND VPWR VPWR _14302_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _15591_/Q VGND VGND VPWR VPWR _12495_/A sky130_fd_sc_hd__inv_2
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15282_ _08610_/X _15282_/D VGND VGND VPWR VPWR _15282_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14233_ _14664_/Q _15240_/Q _14728_/Q _14696_/Q _14265_/S0 _14265_/S1 VGND VGND VPWR
+ VPWR _14233_/X sky130_fd_sc_hd__mux4_2
X_11445_ _11454_/A VGND VGND VPWR VPWR _11445_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14164_ _15183_/Q _15151_/Q _14767_/Q _14799_/Q _14180_/S0 _14210_/S1 VGND VGND VPWR
+ VPWR _14164_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11376_ _14579_/Q _11374_/X _11134_/X _11375_/X VGND VGND VPWR VPWR _14579_/D sky130_fd_sc_hd__a22o_1
X_13115_ _15661_/Q data_address[26] _15667_/Q VGND VGND VPWR VPWR _13115_/X sky130_fd_sc_hd__mux2_1
X_10327_ _10339_/A VGND VGND VPWR VPWR _10327_/X sky130_fd_sc_hd__buf_1
XFILLER_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14095_ _15126_/Q _15350_/Q _15318_/Q _15286_/Q _14145_/S0 _14238_/S1 VGND VGND VPWR
+ VPWR _14095_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13046_ wdata[19] rdata[19] _13058_/S VGND VGND VPWR VPWR _14323_/D sky130_fd_sc_hd__mux2_1
X_10258_ _10258_/A VGND VGND VPWR VPWR _10281_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10189_ _10193_/A VGND VGND VPWR VPWR _10189_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14997_ _09750_/X _14997_/D VGND VGND VPWR VPWR _14997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13948_ _14501_/Q _14469_/Q _14437_/Q _14405_/Q _13950_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13948_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13879_ _14828_/Q _14860_/Q _14892_/Q _14924_/Q _13919_/S0 _13950_/S1 VGND VGND VPWR
+ VPWR _13879_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15618_ _15647_/CLK _15618_/D VGND VGND VPWR VPWR pc[13] sky130_fd_sc_hd__dfxtp_2
XFILLER_148_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15549_ _15592_/CLK _15549_/D VGND VGND VPWR VPWR _15549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09070_ _09074_/A VGND VGND VPWR VPWR _09070_/X sky130_fd_sc_hd__clkbuf_1
X_08021_ _08021_/A VGND VGND VPWR VPWR _08021_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09972_ _09972_/A VGND VGND VPWR VPWR _09972_/X sky130_fd_sc_hd__buf_1
XFILLER_39_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08923_ _08923_/A VGND VGND VPWR VPWR _11062_/B sky130_fd_sc_hd__buf_1
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08854_ _15219_/Q _08851_/X _08852_/X _08853_/X VGND VGND VPWR VPWR _15219_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07805_ _07805_/A _07805_/B VGND VGND VPWR VPWR _07805_/Y sky130_fd_sc_hd__nand2_1
X_08785_ _08800_/A VGND VGND VPWR VPWR _08786_/A sky130_fd_sc_hd__buf_1
XFILLER_84_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07736_ _13144_/X _07730_/B _07731_/A VGND VGND VPWR VPWR _07875_/A sky130_fd_sc_hd__a21oi_1
XFILLER_44_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07667_ _07663_/X _13123_/X _07663_/A _13123_/X VGND VGND VPWR VPWR _07668_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09406_ _15075_/Q _09298_/A _09290_/X _09301_/A VGND VGND VPWR VPWR _15075_/D sky130_fd_sc_hd__a22o_1
X_07598_ _07599_/A _13069_/X VGND VGND VPWR VPWR _15484_/D sky130_fd_sc_hd__and2_1
XFILLER_25_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09337_ _15097_/Q _09335_/X _09196_/X _09336_/X VGND VGND VPWR VPWR _15097_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09268_ _15113_/Q _09262_/X _09267_/X _09264_/X VGND VGND VPWR VPWR _15113_/D sky130_fd_sc_hd__a22o_1
X_08219_ _14301_/Q VGND VGND VPWR VPWR _08662_/C sky130_fd_sc_hd__inv_2
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09199_ _09199_/A VGND VGND VPWR VPWR _09199_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11230_ _11239_/A VGND VGND VPWR VPWR _11237_/A sky130_fd_sc_hd__buf_1
XFILLER_153_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11161_ _11528_/A VGND VGND VPWR VPWR _11161_/X sky130_fd_sc_hd__buf_1
XFILLER_122_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10112_ _14903_/Q _10106_/X _09981_/X _10107_/X VGND VGND VPWR VPWR _14903_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11092_ _14653_/Q _11080_/X _11091_/X _11084_/X VGND VGND VPWR VPWR _14653_/D sky130_fd_sc_hd__a22o_1
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14920_ _10046_/X _14920_/D VGND VGND VPWR VPWR _14920_/Q sky130_fd_sc_hd__dfxtp_1
X_10043_ _14921_/Q _10037_/X _10042_/X _10039_/X VGND VGND VPWR VPWR _14921_/D sky130_fd_sc_hd__a22o_1
XFILLER_121_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14851_ _10291_/X _14851_/D VGND VGND VPWR VPWR _14851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13802_ _15219_/Q _14547_/Q _14995_/Q _15411_/Q _13825_/S0 _13918_/S1 VGND VGND VPWR
+ VPWR _13802_/X sky130_fd_sc_hd__mux4_2
XFILLER_91_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14782_ _10570_/X _14782_/D VGND VGND VPWR VPWR _14782_/Q sky130_fd_sc_hd__dfxtp_1
X_11994_ _11994_/A VGND VGND VPWR VPWR _12001_/A sky130_fd_sc_hd__buf_1
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13733_ _14682_/Q _15258_/Q _14746_/Q _14714_/Q _13737_/S0 _13963_/S1 VGND VGND VPWR
+ VPWR _13733_/X sky130_fd_sc_hd__mux4_2
XFILLER_17_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10945_ _14692_/Q _10840_/A _10828_/X _10843_/A VGND VGND VPWR VPWR _14692_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13664_ _15201_/Q _15169_/Q _14785_/Q _14817_/Q _13740_/S0 _07541_/A VGND VGND VPWR
+ VPWR _13664_/X sky130_fd_sc_hd__mux4_2
X_10876_ _14713_/Q _10874_/X _10718_/X _10875_/X VGND VGND VPWR VPWR _14713_/D sky130_fd_sc_hd__a22o_1
X_15403_ _08057_/X _15403_/D VGND VGND VPWR VPWR _15403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12615_ _15550_/Q VGND VGND VPWR VPWR _12615_/X sky130_fd_sc_hd__buf_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ _13594_/X _13073_/X _14337_/Q VGND VGND VPWR VPWR _13595_/X sky130_fd_sc_hd__mux2_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15334_ _08330_/X _15334_/D VGND VGND VPWR VPWR _15334_/Q sky130_fd_sc_hd__dfxtp_1
X_12546_ _12546_/A VGND VGND VPWR VPWR _12546_/X sky130_fd_sc_hd__buf_1
XFILLER_12_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15265_ _08672_/X _15265_/D VGND VGND VPWR VPWR _15265_/Q sky130_fd_sc_hd__dfxtp_1
X_12477_ _12463_/X _12470_/X _12472_/X _12476_/X VGND VGND VPWR VPWR _12477_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_144_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_4 data_address[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14216_ _14212_/X _14213_/X _14214_/X _14215_/X _14266_/S0 _14266_/S1 VGND VGND VPWR
+ VPWR _14216_/X sky130_fd_sc_hd__mux4_2
X_11428_ _11428_/A _11428_/B VGND VGND VPWR VPWR _11446_/A sky130_fd_sc_hd__or2_2
X_15196_ _08953_/X _15196_/D VGND VGND VPWR VPWR _15196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_14147_ _14641_/Q _14609_/Q _14577_/Q _15377_/Q _14180_/S0 _14396_/Q VGND VGND VPWR
+ VPWR _14147_/X sky130_fd_sc_hd__mux4_1
X_11359_ _14584_/Q _11354_/X _11112_/X _11355_/X VGND VGND VPWR VPWR _14584_/D sky130_fd_sc_hd__a22o_1
XFILLER_112_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14078_ _14520_/Q _14488_/Q _14456_/Q _14424_/Q _14283_/S0 _14284_/S1 VGND VGND VPWR
+ VPWR _14078_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13029_ wdata[2] rdata[2] _13058_/S VGND VGND VPWR VPWR _14306_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08570_ _08572_/A VGND VGND VPWR VPWR _08570_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07521_ _07521_/A VGND VGND VPWR VPWR _07641_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07452_ _07456_/A VGND VGND VPWR VPWR _07455_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07383_ _07383_/A VGND VGND VPWR VPWR _07496_/A sky130_fd_sc_hd__buf_1
XFILLER_50_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09122_ _15148_/Q _09116_/X _08883_/X _09118_/X VGND VGND VPWR VPWR _15148_/D sky130_fd_sc_hd__a22o_1
XFILLER_31_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09053_ _09115_/A VGND VGND VPWR VPWR _09075_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08004_ _08004_/A VGND VGND VPWR VPWR _08004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09955_ _14941_/Q _09943_/X _09954_/X _09947_/X VGND VGND VPWR VPWR _14941_/D sky130_fd_sc_hd__a22o_1
XFILLER_103_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08906_ _08906_/A VGND VGND VPWR VPWR _08906_/X sky130_fd_sc_hd__buf_1
XFILLER_58_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09886_ _09886_/A VGND VGND VPWR VPWR _09907_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08837_ _08876_/A VGND VGND VPWR VPWR _08864_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08768_ _08770_/A VGND VGND VPWR VPWR _08768_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07719_ _13141_/X VGND VGND VPWR VPWR _07720_/A sky130_fd_sc_hd__inv_2
X_08699_ _08701_/A VGND VGND VPWR VPWR _08699_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10730_ _10738_/A VGND VGND VPWR VPWR _10730_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10661_ _11798_/A _10949_/A VGND VGND VPWR VPWR _10680_/A sky130_fd_sc_hd__or2_2
X_12400_ _13329_/X _12400_/B VGND VGND VPWR VPWR _12400_/X sky130_fd_sc_hd__or2_2
X_13380_ _12758_/A _12737_/A _13418_/S VGND VGND VPWR VPWR _13380_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10592_ _14776_/Q _10584_/X _10344_/X _10585_/X VGND VGND VPWR VPWR _14776_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12331_ _12020_/X _12021_/X _12329_/X _12330_/X VGND VGND VPWR VPWR _12904_/A sky130_fd_sc_hd__o22a_1
XFILLER_127_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12262_ _12837_/A _12261_/A _12854_/A _12261_/Y VGND VGND VPWR VPWR _12799_/A sky130_fd_sc_hd__o22a_1
X_15050_ _09495_/X _15050_/D VGND VGND VPWR VPWR _15050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14001_ _13997_/X _13998_/X _13999_/X _14000_/X _14397_/Q _14398_/Q VGND VGND VPWR
+ VPWR _14001_/X sky130_fd_sc_hd__mux4_1
X_11213_ _14625_/Q _11207_/X _11071_/X _11210_/X VGND VGND VPWR VPWR _14625_/D sky130_fd_sc_hd__a22o_1
X_12193_ _12193_/A _12749_/A VGND VGND VPWR VPWR _12209_/A sky130_fd_sc_hd__nand2_1
XFILLER_122_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11144_ _11510_/A VGND VGND VPWR VPWR _11144_/X sky130_fd_sc_hd__buf_1
XFILLER_150_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11075_ _11443_/A VGND VGND VPWR VPWR _11075_/X sky130_fd_sc_hd__buf_1
XFILLER_95_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10026_ _10026_/A VGND VGND VPWR VPWR _10052_/A sky130_fd_sc_hd__clkbuf_2
X_14903_ _10111_/X _14903_/D VGND VGND VPWR VPWR _14903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14834_ _10370_/X _14834_/D VGND VGND VPWR VPWR _14834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14765_ _10625_/X _14765_/D VGND VGND VPWR VPWR _14765_/Q sky130_fd_sc_hd__dfxtp_1
X_11977_ _11977_/A VGND VGND VPWR VPWR _11977_/X sky130_fd_sc_hd__buf_1
XFILLER_72_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13716_ _13712_/X _13713_/X _13714_/X _13715_/X _13966_/S0 _13966_/S1 VGND VGND VPWR
+ VPWR _13716_/X sky130_fd_sc_hd__mux4_2
X_10928_ _14697_/Q _10924_/X _10804_/X _10925_/X VGND VGND VPWR VPWR _14697_/D sky130_fd_sc_hd__a22o_1
X_14696_ _10929_/X _14696_/D VGND VGND VPWR VPWR _14696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13647_ _13646_/X _13060_/X _14337_/Q VGND VGND VPWR VPWR _13647_/X sky130_fd_sc_hd__mux2_1
X_10859_ _14718_/Q _10853_/X _10691_/X _10856_/X VGND VGND VPWR VPWR _14718_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13578_ _13577_/X _14322_/D _15506_/Q VGND VGND VPWR VPWR _13578_/X sky130_fd_sc_hd__mux2_1
X_15317_ _08431_/X _15317_/D VGND VGND VPWR VPWR _15317_/Q sky130_fd_sc_hd__dfxtp_1
X_12529_ _12492_/A _12507_/A _12513_/Y VGND VGND VPWR VPWR _12530_/A sky130_fd_sc_hd__o21ai_2
XFILLER_117_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15248_ _08731_/X _15248_/D VGND VGND VPWR VPWR _15248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15179_ _09012_/X _15179_/D VGND VGND VPWR VPWR _15179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09740_ _15000_/Q _09736_/X _09584_/X _09737_/X VGND VGND VPWR VPWR _15000_/D sky130_fd_sc_hd__a22o_1
.ends

