module core (clk,
    ren,
    rst,
    wen,
    VPWR,
    VGND,
    data_address,
    instruction,
    pc,
    rdata,
    wdata,
    wstrobe);
 input clk;
 output ren;
 input rst;
 output wen;
 input VPWR;
 input VGND;
 output [31:0] data_address;
 input [31:0] instruction;
 output [31:0] pc;
 input [31:0] rdata;
 output [31:0] wdata;
 output [3:0] wstrobe;

 sky130_fd_sc_hd__buf_1 _07105_ (.A(MEM_X_BRANCH_TAKEN),
    .X(_03664_));
 sky130_fd_sc_hd__buf_1 _07106_ (.A(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__inv_2 _07107_ (.A(MEM_X_BRANCH_TAKEN),
    .Y(_03666_));
 sky130_fd_sc_hd__buf_1 _07108_ (.A(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__buf_1 _07109_ (.A(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__buf_1 _07110_ (.A(_03668_),
    .X(_03669_));
 sky130_fd_sc_hd__inv_2 _07111_ (.A(rst),
    .Y(_03670_));
 sky130_fd_sc_hd__clkbuf_2 _07112_ (.A(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__buf_1 _07113_ (.A(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__o221a_1 _07114_ (.A1(_03665_),
    .A2(\next_pc[0] ),
    .B1(_03669_),
    .B2(data_address[0]),
    .C1(_03672_),
    .X(_03662_));
 sky130_fd_sc_hd__clkbuf_1 _07115_ (.A(_03667_),
    .X(_03673_));
 sky130_fd_sc_hd__buf_1 _07116_ (.A(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__buf_1 _07117_ (.A(\c1.instruction2[6] ),
    .X(_03675_));
 sky130_fd_sc_hd__inv_2 _07118_ (.A(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__inv_2 _07119_ (.A(\c1.instruction2[5] ),
    .Y(_03677_));
 sky130_fd_sc_hd__or4bb_4 _07120_ (.A(\c1.instruction2[3] ),
    .B(\c1.instruction2[2] ),
    .C_N(\c1.instruction2[1] ),
    .D_N(\c1.instruction2[0] ),
    .X(_03678_));
 sky130_fd_sc_hd__buf_1 _07121_ (.A(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__or4_4 _07122_ (.A(_03676_),
    .B(_03677_),
    .C(\c1.instruction2[4] ),
    .D(_03679_),
    .X(_03680_));
 sky130_fd_sc_hd__inv_16 _07123_ (.A(_03680_),
    .Y(_00014_));
 sky130_fd_sc_hd__and3_1 _07124_ (.A(_03674_),
    .B(\e1.alu1.out[0] ),
    .C(_00014_),
    .X(_03661_));
 sky130_fd_sc_hd__inv_2 _07125_ (.A(_01359_),
    .Y(_03681_));
 sky130_fd_sc_hd__inv_2 _07126_ (.A(_01358_),
    .Y(_03682_));
 sky130_fd_sc_hd__inv_2 _07127_ (.A(_01357_),
    .Y(_03683_));
 sky130_fd_sc_hd__inv_2 _07128_ (.A(_01356_),
    .Y(_03684_));
 sky130_fd_sc_hd__inv_2 _07129_ (.A(_01355_),
    .Y(_03685_));
 sky130_fd_sc_hd__inv_2 _07130_ (.A(_01354_),
    .Y(_03686_));
 sky130_fd_sc_hd__inv_2 _07131_ (.A(_01353_),
    .Y(_03687_));
 sky130_fd_sc_hd__inv_2 _07132_ (.A(_01352_),
    .Y(_03688_));
 sky130_fd_sc_hd__inv_2 _07133_ (.A(_01351_),
    .Y(_03689_));
 sky130_fd_sc_hd__inv_2 _07134_ (.A(_01349_),
    .Y(_03690_));
 sky130_fd_sc_hd__inv_2 _07135_ (.A(_01348_),
    .Y(_03691_));
 sky130_fd_sc_hd__inv_2 _07136_ (.A(_01347_),
    .Y(_03692_));
 sky130_fd_sc_hd__inv_2 _07137_ (.A(_01346_),
    .Y(_03693_));
 sky130_fd_sc_hd__inv_2 _07138_ (.A(_01345_),
    .Y(_03694_));
 sky130_fd_sc_hd__inv_2 _07139_ (.A(_01344_),
    .Y(_03695_));
 sky130_fd_sc_hd__inv_2 _07140_ (.A(_01343_),
    .Y(_03696_));
 sky130_fd_sc_hd__inv_2 _07141_ (.A(_01342_),
    .Y(_03697_));
 sky130_fd_sc_hd__inv_2 _07142_ (.A(_01341_),
    .Y(_03698_));
 sky130_fd_sc_hd__inv_2 _07143_ (.A(_01340_),
    .Y(_03699_));
 sky130_fd_sc_hd__inv_2 _07144_ (.A(_01368_),
    .Y(_03700_));
 sky130_fd_sc_hd__inv_2 _07145_ (.A(_01367_),
    .Y(_03701_));
 sky130_fd_sc_hd__inv_2 _07146_ (.A(_01366_),
    .Y(_03702_));
 sky130_fd_sc_hd__inv_2 _07147_ (.A(_01365_),
    .Y(_03703_));
 sky130_fd_sc_hd__inv_2 _07148_ (.A(_01364_),
    .Y(_03704_));
 sky130_fd_sc_hd__inv_2 _07149_ (.A(_01363_),
    .Y(_03705_));
 sky130_fd_sc_hd__inv_2 _07150_ (.A(_01350_),
    .Y(_03706_));
 sky130_fd_sc_hd__inv_2 _07151_ (.A(_01339_),
    .Y(_03707_));
 sky130_fd_sc_hd__inv_2 _07152_ (.A(_01361_),
    .Y(_03708_));
 sky130_fd_sc_hd__inv_2 _07153_ (.A(_01362_),
    .Y(_03709_));
 sky130_fd_sc_hd__or4_4 _07154_ (.A(_03706_),
    .B(_03707_),
    .C(_03708_),
    .D(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__or2_1 _07155_ (.A(_03705_),
    .B(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__or2_2 _07156_ (.A(_03704_),
    .B(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__or2_1 _07157_ (.A(_03703_),
    .B(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__or2_1 _07158_ (.A(_03702_),
    .B(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__or2_1 _07159_ (.A(_03701_),
    .B(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__or2_1 _07160_ (.A(_03700_),
    .B(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__or2_1 _07161_ (.A(_03699_),
    .B(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__or2_2 _07162_ (.A(_03698_),
    .B(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__or2_1 _07163_ (.A(_03697_),
    .B(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__or2_2 _07164_ (.A(_03696_),
    .B(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__or2_1 _07165_ (.A(_03695_),
    .B(_03720_),
    .X(_03721_));
 sky130_fd_sc_hd__or2_2 _07166_ (.A(_03694_),
    .B(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__or2_1 _07167_ (.A(_03693_),
    .B(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__or2_4 _07168_ (.A(_03692_),
    .B(_03723_),
    .X(_03724_));
 sky130_fd_sc_hd__or2_1 _07169_ (.A(_03691_),
    .B(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__or2_1 _07170_ (.A(_03690_),
    .B(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__or2_1 _07171_ (.A(_03689_),
    .B(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__or2_2 _07172_ (.A(_03688_),
    .B(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__or2_1 _07173_ (.A(_03687_),
    .B(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__or2_2 _07174_ (.A(_03686_),
    .B(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__or2_1 _07175_ (.A(_03685_),
    .B(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__or2_2 _07176_ (.A(_03684_),
    .B(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__or2_1 _07177_ (.A(_03683_),
    .B(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__or2_2 _07178_ (.A(_03682_),
    .B(_03733_),
    .X(_03734_));
 sky130_fd_sc_hd__or2_1 _07179_ (.A(_03681_),
    .B(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__inv_2 _07180_ (.A(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__inv_2 _07181_ (.A(_01360_),
    .Y(_03737_));
 sky130_fd_sc_hd__buf_1 _07182_ (.A(_03670_),
    .X(_03738_));
 sky130_fd_sc_hd__buf_1 _07183_ (.A(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__buf_1 _07184_ (.A(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__o221a_1 _07185_ (.A1(_01360_),
    .A2(_03736_),
    .B1(_03737_),
    .B2(_03735_),
    .C1(_03740_),
    .X(_03660_));
 sky130_fd_sc_hd__buf_1 _07186_ (.A(rst),
    .X(_03741_));
 sky130_fd_sc_hd__buf_1 _07187_ (.A(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__buf_2 _07188_ (.A(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__a211oi_2 _07189_ (.A1(_03681_),
    .A2(_03734_),
    .B1(_03743_),
    .C1(_03736_),
    .Y(_03659_));
 sky130_fd_sc_hd__inv_2 _07190_ (.A(_03733_),
    .Y(_03744_));
 sky130_fd_sc_hd__buf_1 _07191_ (.A(_03738_),
    .X(_03745_));
 sky130_fd_sc_hd__o211a_1 _07192_ (.A1(_01358_),
    .A2(_03744_),
    .B1(_03745_),
    .C1(_03734_),
    .X(_03658_));
 sky130_fd_sc_hd__a211oi_2 _07193_ (.A1(_03683_),
    .A2(_03732_),
    .B1(_03743_),
    .C1(_03744_),
    .Y(_03657_));
 sky130_fd_sc_hd__inv_2 _07194_ (.A(_03731_),
    .Y(_03746_));
 sky130_fd_sc_hd__o211a_1 _07195_ (.A1(_01356_),
    .A2(_03746_),
    .B1(_03745_),
    .C1(_03732_),
    .X(_03656_));
 sky130_fd_sc_hd__a211oi_4 _07196_ (.A1(_03685_),
    .A2(_03730_),
    .B1(_03743_),
    .C1(_03746_),
    .Y(_03655_));
 sky130_fd_sc_hd__inv_2 _07197_ (.A(_03729_),
    .Y(_03747_));
 sky130_fd_sc_hd__buf_1 _07198_ (.A(_03671_),
    .X(_03748_));
 sky130_fd_sc_hd__o211a_1 _07199_ (.A1(_01354_),
    .A2(_03747_),
    .B1(_03748_),
    .C1(_03730_),
    .X(_03654_));
 sky130_fd_sc_hd__buf_2 _07200_ (.A(_03742_),
    .X(_03749_));
 sky130_fd_sc_hd__a211oi_4 _07201_ (.A1(_03687_),
    .A2(_03728_),
    .B1(_03749_),
    .C1(_03747_),
    .Y(_03653_));
 sky130_fd_sc_hd__inv_2 _07202_ (.A(_03727_),
    .Y(_03750_));
 sky130_fd_sc_hd__o211a_1 _07203_ (.A1(_01352_),
    .A2(_03750_),
    .B1(_03748_),
    .C1(_03728_),
    .X(_03652_));
 sky130_fd_sc_hd__a211oi_2 _07204_ (.A1(_03689_),
    .A2(_03726_),
    .B1(_03749_),
    .C1(_03750_),
    .Y(_03651_));
 sky130_fd_sc_hd__inv_2 _07205_ (.A(_03725_),
    .Y(_03751_));
 sky130_fd_sc_hd__o211a_1 _07206_ (.A1(_01349_),
    .A2(_03751_),
    .B1(_03748_),
    .C1(_03726_),
    .X(_03650_));
 sky130_fd_sc_hd__a211oi_2 _07207_ (.A1(_03691_),
    .A2(_03724_),
    .B1(_03749_),
    .C1(_03751_),
    .Y(_03649_));
 sky130_fd_sc_hd__inv_2 _07208_ (.A(_03723_),
    .Y(_03752_));
 sky130_fd_sc_hd__buf_1 _07209_ (.A(_03671_),
    .X(_03753_));
 sky130_fd_sc_hd__o211a_1 _07210_ (.A1(_01347_),
    .A2(_03752_),
    .B1(_03753_),
    .C1(_03724_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_1 _07211_ (.A(_03741_),
    .X(_03754_));
 sky130_fd_sc_hd__buf_2 _07212_ (.A(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__a211oi_2 _07213_ (.A1(_03693_),
    .A2(_03722_),
    .B1(_03755_),
    .C1(_03752_),
    .Y(_03647_));
 sky130_fd_sc_hd__inv_2 _07214_ (.A(_03721_),
    .Y(_03756_));
 sky130_fd_sc_hd__o211a_1 _07215_ (.A1(_01345_),
    .A2(_03756_),
    .B1(_03753_),
    .C1(_03722_),
    .X(_03646_));
 sky130_fd_sc_hd__a211oi_2 _07216_ (.A1(_03695_),
    .A2(_03720_),
    .B1(_03755_),
    .C1(_03756_),
    .Y(_03645_));
 sky130_fd_sc_hd__inv_2 _07217_ (.A(_03719_),
    .Y(_03757_));
 sky130_fd_sc_hd__o211a_1 _07218_ (.A1(_01343_),
    .A2(_03757_),
    .B1(_03753_),
    .C1(_03720_),
    .X(_03644_));
 sky130_fd_sc_hd__a211oi_2 _07219_ (.A1(_03697_),
    .A2(_03718_),
    .B1(_03755_),
    .C1(_03757_),
    .Y(_03643_));
 sky130_fd_sc_hd__inv_2 _07220_ (.A(_03717_),
    .Y(_03758_));
 sky130_fd_sc_hd__buf_1 _07221_ (.A(_03738_),
    .X(_03759_));
 sky130_fd_sc_hd__o211a_1 _07222_ (.A1(_01341_),
    .A2(_03758_),
    .B1(_03759_),
    .C1(_03718_),
    .X(_03642_));
 sky130_fd_sc_hd__buf_1 _07223_ (.A(_03754_),
    .X(_03760_));
 sky130_fd_sc_hd__a211oi_1 _07224_ (.A1(_03699_),
    .A2(_03716_),
    .B1(_03760_),
    .C1(_03758_),
    .Y(_03641_));
 sky130_fd_sc_hd__inv_2 _07225_ (.A(_03715_),
    .Y(_03761_));
 sky130_fd_sc_hd__o211a_1 _07226_ (.A1(_01368_),
    .A2(_03761_),
    .B1(_03759_),
    .C1(_03716_),
    .X(_03640_));
 sky130_fd_sc_hd__a211oi_2 _07227_ (.A1(_03701_),
    .A2(_03714_),
    .B1(_03760_),
    .C1(_03761_),
    .Y(_03639_));
 sky130_fd_sc_hd__inv_2 _07228_ (.A(_03713_),
    .Y(_03762_));
 sky130_fd_sc_hd__o211a_1 _07229_ (.A1(_01366_),
    .A2(_03762_),
    .B1(_03759_),
    .C1(_03714_),
    .X(_03638_));
 sky130_fd_sc_hd__a211oi_2 _07230_ (.A1(_03703_),
    .A2(_03712_),
    .B1(_03760_),
    .C1(_03762_),
    .Y(_03637_));
 sky130_fd_sc_hd__inv_2 _07231_ (.A(_03711_),
    .Y(_03763_));
 sky130_fd_sc_hd__o211a_1 _07232_ (.A1(_01364_),
    .A2(_03763_),
    .B1(_03739_),
    .C1(_03712_),
    .X(_03636_));
 sky130_fd_sc_hd__inv_2 _07233_ (.A(_03710_),
    .Y(_03764_));
 sky130_fd_sc_hd__o211a_1 _07234_ (.A1(_01363_),
    .A2(_03764_),
    .B1(_03739_),
    .C1(_03711_),
    .X(_03635_));
 sky130_fd_sc_hd__buf_1 _07235_ (.A(_03742_),
    .X(_03765_));
 sky130_fd_sc_hd__buf_1 _07236_ (.A(_03706_),
    .X(_03766_));
 sky130_fd_sc_hd__buf_1 _07237_ (.A(_03707_),
    .X(_03767_));
 sky130_fd_sc_hd__o31a_1 _07238_ (.A1(_03766_),
    .A2(_03767_),
    .A3(_03708_),
    .B1(_03709_),
    .X(_03768_));
 sky130_fd_sc_hd__nor3_1 _07239_ (.A(_03765_),
    .B(_03764_),
    .C(_03768_),
    .Y(_03634_));
 sky130_fd_sc_hd__buf_1 _07240_ (.A(_03766_),
    .X(_03769_));
 sky130_fd_sc_hd__buf_1 _07241_ (.A(_03767_),
    .X(_03770_));
 sky130_fd_sc_hd__buf_1 _07242_ (.A(_03708_),
    .X(_03771_));
 sky130_fd_sc_hd__o21ai_1 _07243_ (.A1(_03766_),
    .A2(_03770_),
    .B1(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__o311a_1 _07244_ (.A1(_03769_),
    .A2(_03770_),
    .A3(_03771_),
    .B1(_03745_),
    .C1(_03772_),
    .X(_03633_));
 sky130_fd_sc_hd__o221a_1 _07245_ (.A1(_03769_),
    .A2(_03770_),
    .B1(_01350_),
    .B2(_01339_),
    .C1(_03740_),
    .X(_03632_));
 sky130_fd_sc_hd__or2_1 _07246_ (.A(_03754_),
    .B(_03767_),
    .X(_03631_));
 sky130_fd_sc_hd__buf_1 _07247_ (.A(_03741_),
    .X(_03773_));
 sky130_fd_sc_hd__buf_1 _07248_ (.A(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_2 _07249_ (.A(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__nor2_1 _07250_ (.A(_03775_),
    .B(_03737_),
    .Y(_03630_));
 sky130_fd_sc_hd__nor2_4 _07251_ (.A(_03775_),
    .B(_03681_),
    .Y(_03629_));
 sky130_fd_sc_hd__nor2_1 _07252_ (.A(_03775_),
    .B(_03682_),
    .Y(_03628_));
 sky130_fd_sc_hd__buf_1 _07253_ (.A(_03774_),
    .X(_03776_));
 sky130_fd_sc_hd__nor2_1 _07254_ (.A(_03776_),
    .B(_03683_),
    .Y(_03627_));
 sky130_fd_sc_hd__nor2_1 _07255_ (.A(_03776_),
    .B(_03684_),
    .Y(_03626_));
 sky130_fd_sc_hd__nor2_1 _07256_ (.A(_03776_),
    .B(_03685_),
    .Y(_03625_));
 sky130_fd_sc_hd__buf_1 _07257_ (.A(_03774_),
    .X(_03777_));
 sky130_fd_sc_hd__nor2_1 _07258_ (.A(_03777_),
    .B(_03686_),
    .Y(_03624_));
 sky130_fd_sc_hd__nor2_1 _07259_ (.A(_03777_),
    .B(_03687_),
    .Y(_03623_));
 sky130_fd_sc_hd__nor2_1 _07260_ (.A(_03777_),
    .B(_03688_),
    .Y(_03622_));
 sky130_fd_sc_hd__clkbuf_2 _07261_ (.A(_03773_),
    .X(_03778_));
 sky130_fd_sc_hd__clkbuf_2 _07262_ (.A(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__nor2_1 _07263_ (.A(_03779_),
    .B(_03689_),
    .Y(_03621_));
 sky130_fd_sc_hd__nor2_1 _07264_ (.A(_03779_),
    .B(_03690_),
    .Y(_03620_));
 sky130_fd_sc_hd__nor2_4 _07265_ (.A(_03779_),
    .B(_03691_),
    .Y(_03619_));
 sky130_fd_sc_hd__buf_1 _07266_ (.A(_03778_),
    .X(_03780_));
 sky130_fd_sc_hd__nor2_1 _07267_ (.A(_03780_),
    .B(_03692_),
    .Y(_03618_));
 sky130_fd_sc_hd__nor2_1 _07268_ (.A(_03780_),
    .B(_03693_),
    .Y(_03617_));
 sky130_fd_sc_hd__nor2_1 _07269_ (.A(_03780_),
    .B(_03694_),
    .Y(_03616_));
 sky130_fd_sc_hd__buf_1 _07270_ (.A(_03778_),
    .X(_03781_));
 sky130_fd_sc_hd__nor2_1 _07271_ (.A(_03781_),
    .B(_03695_),
    .Y(_03615_));
 sky130_fd_sc_hd__nor2_1 _07272_ (.A(_03781_),
    .B(_03696_),
    .Y(_03614_));
 sky130_fd_sc_hd__nor2_1 _07273_ (.A(_03781_),
    .B(_03697_),
    .Y(_03613_));
 sky130_fd_sc_hd__buf_1 _07274_ (.A(_03773_),
    .X(_03782_));
 sky130_fd_sc_hd__buf_1 _07275_ (.A(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__nor2_1 _07276_ (.A(_03783_),
    .B(_03698_),
    .Y(_03612_));
 sky130_fd_sc_hd__nor2_1 _07277_ (.A(_03783_),
    .B(_03699_),
    .Y(_03611_));
 sky130_fd_sc_hd__nor2_1 _07278_ (.A(_03783_),
    .B(_03700_),
    .Y(_03610_));
 sky130_fd_sc_hd__buf_1 _07279_ (.A(_03782_),
    .X(_03784_));
 sky130_fd_sc_hd__nor2_1 _07280_ (.A(_03784_),
    .B(_03701_),
    .Y(_03609_));
 sky130_fd_sc_hd__nor2_1 _07281_ (.A(_03784_),
    .B(_03702_),
    .Y(_03608_));
 sky130_fd_sc_hd__nor2_1 _07282_ (.A(_03784_),
    .B(_03703_),
    .Y(_03607_));
 sky130_fd_sc_hd__buf_1 _07283_ (.A(_03782_),
    .X(_03785_));
 sky130_fd_sc_hd__nor2_1 _07284_ (.A(_03785_),
    .B(_03704_),
    .Y(_03606_));
 sky130_fd_sc_hd__nor2_1 _07285_ (.A(_03785_),
    .B(_03705_),
    .Y(_03605_));
 sky130_fd_sc_hd__nor2_1 _07286_ (.A(_03785_),
    .B(_03709_),
    .Y(_03604_));
 sky130_fd_sc_hd__nor2_1 _07287_ (.A(_03765_),
    .B(_03771_),
    .Y(_03603_));
 sky130_fd_sc_hd__nor2_1 _07288_ (.A(_03765_),
    .B(_03769_),
    .Y(_03602_));
 sky130_fd_sc_hd__inv_2 _07289_ (.A(_03631_),
    .Y(_03601_));
 sky130_fd_sc_hd__and2_1 _07290_ (.A(_03672_),
    .B(_01338_),
    .X(_03600_));
 sky130_fd_sc_hd__and2_1 _07291_ (.A(_03672_),
    .B(_01337_),
    .X(_03599_));
 sky130_fd_sc_hd__inv_2 _07292_ (.A(\c1.instruction1[31] ),
    .Y(_03786_));
 sky130_fd_sc_hd__buf_1 _07293_ (.A(\c1.instruction1[6] ),
    .X(_03787_));
 sky130_fd_sc_hd__inv_2 _07294_ (.A(\c1.instruction1[4] ),
    .Y(_03788_));
 sky130_fd_sc_hd__or4bb_4 _07295_ (.A(\c1.instruction1[3] ),
    .B(\c1.instruction1[2] ),
    .C_N(\c1.instruction1[1] ),
    .D_N(\c1.instruction1[0] ),
    .X(_03789_));
 sky130_fd_sc_hd__or4_4 _07296_ (.A(_03787_),
    .B(\c1.instruction1[5] ),
    .C(_03788_),
    .D(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__buf_1 _07297_ (.A(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__clkbuf_2 _07298_ (.A(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__inv_2 _07299_ (.A(\c1.instruction1[12] ),
    .Y(_03793_));
 sky130_fd_sc_hd__nor2_1 _07300_ (.A(\c1.instruction1[13] ),
    .B(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__clkbuf_2 _07301_ (.A(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__inv_2 _07302_ (.A(\c1.instruction1[5] ),
    .Y(_03796_));
 sky130_fd_sc_hd__buf_1 _07303_ (.A(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__or2_1 _07304_ (.A(\c1.instruction1[4] ),
    .B(_03789_),
    .X(_03798_));
 sky130_fd_sc_hd__clkbuf_1 _07305_ (.A(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__or3_1 _07306_ (.A(\c1.instruction1[6] ),
    .B(\c1.instruction1[5] ),
    .C(_03798_),
    .X(_03800_));
 sky130_fd_sc_hd__buf_1 _07307_ (.A(_03800_),
    .X(_03801_));
 sky130_fd_sc_hd__buf_1 _07308_ (.A(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__o221a_2 _07309_ (.A1(_03792_),
    .A2(_03795_),
    .B1(_03797_),
    .B2(_03799_),
    .C1(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__nor2_8 _07310_ (.A(_03786_),
    .B(_03803_),
    .Y(\d1.addr[11] ));
 sky130_fd_sc_hd__buf_1 _07311_ (.A(MEM_X_BRANCH_TAKEN),
    .X(_03804_));
 sky130_fd_sc_hd__buf_1 _07312_ (.A(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__nor2_1 _07313_ (.A(_03805_),
    .B(_03786_),
    .Y(_03522_));
 sky130_fd_sc_hd__nor2b_1 _07314_ (.A(_03803_),
    .B_N(_03522_),
    .Y(_03598_));
 sky130_fd_sc_hd__inv_2 _07315_ (.A(\c1.instruction1[7] ),
    .Y(_03806_));
 sky130_fd_sc_hd__inv_2 _07316_ (.A(\c1.instruction1[6] ),
    .Y(_03807_));
 sky130_fd_sc_hd__or3_1 _07317_ (.A(_03796_),
    .B(_03799_),
    .C(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__buf_1 _07318_ (.A(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__buf_1 _07319_ (.A(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__inv_2 _07320_ (.A(\c1.instruction1[30] ),
    .Y(_03811_));
 sky130_fd_sc_hd__or3_1 _07321_ (.A(_03787_),
    .B(_03796_),
    .C(_03799_),
    .X(_03812_));
 sky130_fd_sc_hd__buf_1 _07322_ (.A(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__o211a_1 _07323_ (.A1(_03790_),
    .A2(_03794_),
    .B1(_03800_),
    .C1(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__buf_1 _07324_ (.A(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__o22a_1 _07325_ (.A1(_03806_),
    .A2(_03810_),
    .B1(_03811_),
    .B2(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__inv_2 _07326_ (.A(_03816_),
    .Y(\d1.addr[10] ));
 sky130_fd_sc_hd__buf_1 _07327_ (.A(_03664_),
    .X(_03817_));
 sky130_fd_sc_hd__buf_1 _07328_ (.A(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__nor2_1 _07329_ (.A(_03818_),
    .B(_03816_),
    .Y(_03597_));
 sky130_fd_sc_hd__inv_2 _07330_ (.A(\c1.instruction1[29] ),
    .Y(_03819_));
 sky130_fd_sc_hd__o22a_1 _07331_ (.A1(_03811_),
    .A2(_03810_),
    .B1(_03819_),
    .B2(_03815_),
    .X(_03820_));
 sky130_fd_sc_hd__inv_2 _07332_ (.A(_03820_),
    .Y(\d1.addr[9] ));
 sky130_fd_sc_hd__nor2_1 _07333_ (.A(_03818_),
    .B(_03820_),
    .Y(_03596_));
 sky130_fd_sc_hd__inv_2 _07334_ (.A(\c1.instruction1[28] ),
    .Y(_03821_));
 sky130_fd_sc_hd__o22a_1 _07335_ (.A1(_03819_),
    .A2(_03810_),
    .B1(_03821_),
    .B2(_03815_),
    .X(_03822_));
 sky130_fd_sc_hd__inv_2 _07336_ (.A(_03822_),
    .Y(\d1.addr[8] ));
 sky130_fd_sc_hd__nor2_1 _07337_ (.A(_03818_),
    .B(_03822_),
    .Y(_03595_));
 sky130_fd_sc_hd__buf_1 _07338_ (.A(_03808_),
    .X(_03823_));
 sky130_fd_sc_hd__buf_1 _07339_ (.A(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__inv_2 _07340_ (.A(\c1.instruction1[27] ),
    .Y(_03825_));
 sky130_fd_sc_hd__buf_1 _07341_ (.A(_03814_),
    .X(_03826_));
 sky130_fd_sc_hd__o22a_1 _07342_ (.A1(_03821_),
    .A2(_03824_),
    .B1(_03825_),
    .B2(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__inv_2 _07343_ (.A(_03827_),
    .Y(\d1.addr[7] ));
 sky130_fd_sc_hd__buf_1 _07344_ (.A(_03817_),
    .X(_03828_));
 sky130_fd_sc_hd__nor2_1 _07345_ (.A(_03828_),
    .B(_03827_),
    .Y(_03594_));
 sky130_fd_sc_hd__inv_2 _07346_ (.A(\c1.instruction1[26] ),
    .Y(_03829_));
 sky130_fd_sc_hd__o22a_1 _07347_ (.A1(_03825_),
    .A2(_03824_),
    .B1(_03829_),
    .B2(_03826_),
    .X(_03830_));
 sky130_fd_sc_hd__inv_2 _07348_ (.A(_03830_),
    .Y(\d1.addr[6] ));
 sky130_fd_sc_hd__nor2_1 _07349_ (.A(_03828_),
    .B(_03830_),
    .Y(_03593_));
 sky130_fd_sc_hd__inv_2 _07350_ (.A(\c1.instruction1[25] ),
    .Y(_03831_));
 sky130_fd_sc_hd__o22a_2 _07351_ (.A1(_03829_),
    .A2(_03824_),
    .B1(_03831_),
    .B2(_03826_),
    .X(_03832_));
 sky130_fd_sc_hd__inv_2 _07352_ (.A(_03832_),
    .Y(\d1.addr[5] ));
 sky130_fd_sc_hd__nor2_1 _07353_ (.A(_03828_),
    .B(_03832_),
    .Y(_03592_));
 sky130_fd_sc_hd__buf_1 _07354_ (.A(_03823_),
    .X(_03833_));
 sky130_fd_sc_hd__inv_2 _07355_ (.A(\c1.instruction1[11] ),
    .Y(_03834_));
 sky130_fd_sc_hd__buf_1 _07356_ (.A(_03812_),
    .X(_03835_));
 sky130_fd_sc_hd__inv_2 _07357_ (.A(net53),
    .Y(_03836_));
 sky130_fd_sc_hd__o22a_1 _07358_ (.A1(_03834_),
    .A2(_03835_),
    .B1(_03836_),
    .B2(_03802_),
    .X(_03837_));
 sky130_fd_sc_hd__o221a_2 _07359_ (.A1(_00408_),
    .A2(_03792_),
    .B1(_03831_),
    .B2(_03833_),
    .C1(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__inv_2 _07360_ (.A(_03838_),
    .Y(\d1.addr[4] ));
 sky130_fd_sc_hd__buf_1 _07361_ (.A(_03817_),
    .X(_03839_));
 sky130_fd_sc_hd__nor2_1 _07362_ (.A(_03839_),
    .B(_03838_),
    .Y(_03591_));
 sky130_fd_sc_hd__buf_1 _07363_ (.A(_03791_),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _07364_ (.A(\c1.instruction1[10] ),
    .Y(_03841_));
 sky130_fd_sc_hd__inv_2 _07365_ (.A(\c1.instruction1[23] ),
    .Y(_03842_));
 sky130_fd_sc_hd__buf_1 _07366_ (.A(_03842_),
    .X(_00403_));
 sky130_fd_sc_hd__o22a_1 _07367_ (.A1(_03841_),
    .A2(_03835_),
    .B1(_00403_),
    .B2(_03802_),
    .X(_03843_));
 sky130_fd_sc_hd__o221a_2 _07368_ (.A1(_00405_),
    .A2(_03840_),
    .B1(_03834_),
    .B2(_03833_),
    .C1(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__inv_2 _07369_ (.A(_03844_),
    .Y(\d1.addr[3] ));
 sky130_fd_sc_hd__nor2_1 _07370_ (.A(_03839_),
    .B(_03844_),
    .Y(_03590_));
 sky130_fd_sc_hd__inv_2 _07371_ (.A(\c1.instruction1[9] ),
    .Y(_03845_));
 sky130_fd_sc_hd__inv_2 _07372_ (.A(\c1.instruction1[22] ),
    .Y(_03846_));
 sky130_fd_sc_hd__buf_1 _07373_ (.A(_03801_),
    .X(_03847_));
 sky130_fd_sc_hd__o22a_1 _07374_ (.A1(_03845_),
    .A2(_03835_),
    .B1(_03846_),
    .B2(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__o221a_2 _07375_ (.A1(_00402_),
    .A2(_03840_),
    .B1(_03841_),
    .B2(_03833_),
    .C1(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__inv_2 _07376_ (.A(_03849_),
    .Y(\d1.addr[2] ));
 sky130_fd_sc_hd__nor2_1 _07377_ (.A(_03839_),
    .B(_03849_),
    .Y(_03589_));
 sky130_fd_sc_hd__inv_2 _07378_ (.A(\c1.instruction1[8] ),
    .Y(_03850_));
 sky130_fd_sc_hd__inv_2 _07379_ (.A(net40),
    .Y(_03851_));
 sky130_fd_sc_hd__o22a_1 _07380_ (.A1(_03850_),
    .A2(_03813_),
    .B1(_03851_),
    .B2(_03847_),
    .X(_03852_));
 sky130_fd_sc_hd__o221a_2 _07381_ (.A1(_00399_),
    .A2(_03840_),
    .B1(_03845_),
    .B2(_03809_),
    .C1(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__inv_2 _07382_ (.A(_03853_),
    .Y(\d1.addr[1] ));
 sky130_fd_sc_hd__buf_1 _07383_ (.A(_03664_),
    .X(_03854_));
 sky130_fd_sc_hd__buf_1 _07384_ (.A(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__nor2_1 _07385_ (.A(_03855_),
    .B(_03853_),
    .Y(_03588_));
 sky130_fd_sc_hd__inv_2 _07386_ (.A(_00396_),
    .Y(_03856_));
 sky130_fd_sc_hd__inv_2 _07387_ (.A(net50),
    .Y(_03857_));
 sky130_fd_sc_hd__buf_1 _07388_ (.A(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__o22a_1 _07389_ (.A1(_03806_),
    .A2(_03813_),
    .B1(_03858_),
    .B2(_03847_),
    .X(_03859_));
 sky130_fd_sc_hd__o221a_2 _07390_ (.A1(_03856_),
    .A2(_03791_),
    .B1(_03850_),
    .B2(_03809_),
    .C1(_03859_),
    .X(_03860_));
 sky130_fd_sc_hd__inv_2 _07391_ (.A(_03860_),
    .Y(\d1.addr[0] ));
 sky130_fd_sc_hd__nor2_1 _07392_ (.A(_03855_),
    .B(_03860_),
    .Y(_03587_));
 sky130_fd_sc_hd__buf_1 _07393_ (.A(_03666_),
    .X(_03861_));
 sky130_fd_sc_hd__buf_1 _07394_ (.A(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__clkbuf_2 _07395_ (.A(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__buf_1 _07396_ (.A(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__and2_1 _07397_ (.A(_03864_),
    .B(_01297_),
    .X(_03586_));
 sky130_fd_sc_hd__and2_1 _07398_ (.A(_03864_),
    .B(_01296_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_1 _07399_ (.A(_03863_),
    .X(_03865_));
 sky130_fd_sc_hd__and2_1 _07400_ (.A(_03865_),
    .B(_01294_),
    .X(_03584_));
 sky130_fd_sc_hd__and2_1 _07401_ (.A(_03865_),
    .B(_01293_),
    .X(_03583_));
 sky130_fd_sc_hd__and2_1 _07402_ (.A(_03865_),
    .B(_01292_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_1 _07403_ (.A(_03863_),
    .X(_03866_));
 sky130_fd_sc_hd__and2_1 _07404_ (.A(_03866_),
    .B(_01291_),
    .X(_03581_));
 sky130_fd_sc_hd__and2_1 _07405_ (.A(_03866_),
    .B(_01290_),
    .X(_03580_));
 sky130_fd_sc_hd__and2_1 _07406_ (.A(_03866_),
    .B(_01289_),
    .X(_03579_));
 sky130_fd_sc_hd__clkbuf_2 _07407_ (.A(_03862_),
    .X(_03867_));
 sky130_fd_sc_hd__buf_1 _07408_ (.A(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__and2_1 _07409_ (.A(_03868_),
    .B(_01288_),
    .X(_03578_));
 sky130_fd_sc_hd__and2_1 _07410_ (.A(_03868_),
    .B(_01287_),
    .X(_03577_));
 sky130_fd_sc_hd__and2_1 _07411_ (.A(_03868_),
    .B(_01286_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_1 _07412_ (.A(_03867_),
    .X(_03869_));
 sky130_fd_sc_hd__and2_1 _07413_ (.A(_03869_),
    .B(_01285_),
    .X(_03575_));
 sky130_fd_sc_hd__and2_1 _07414_ (.A(_03869_),
    .B(_01283_),
    .X(_03574_));
 sky130_fd_sc_hd__and2_1 _07415_ (.A(_03869_),
    .B(_01282_),
    .X(_03573_));
 sky130_fd_sc_hd__buf_1 _07416_ (.A(_03867_),
    .X(_03870_));
 sky130_fd_sc_hd__and2_1 _07417_ (.A(_03870_),
    .B(_01281_),
    .X(_03572_));
 sky130_fd_sc_hd__and2_1 _07418_ (.A(_03870_),
    .B(_01280_),
    .X(_03571_));
 sky130_fd_sc_hd__and2_1 _07419_ (.A(_03870_),
    .B(_01279_),
    .X(_03570_));
 sky130_fd_sc_hd__buf_1 _07420_ (.A(_03862_),
    .X(_03871_));
 sky130_fd_sc_hd__clkbuf_1 _07421_ (.A(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__and2_1 _07422_ (.A(_03872_),
    .B(_01278_),
    .X(_03569_));
 sky130_fd_sc_hd__and2_1 _07423_ (.A(_03872_),
    .B(_01277_),
    .X(_03568_));
 sky130_fd_sc_hd__and2_1 _07424_ (.A(_03872_),
    .B(_01276_),
    .X(_03567_));
 sky130_fd_sc_hd__clkbuf_1 _07425_ (.A(_03871_),
    .X(_03873_));
 sky130_fd_sc_hd__and2_1 _07426_ (.A(_03873_),
    .B(_01275_),
    .X(_03566_));
 sky130_fd_sc_hd__and2_1 _07427_ (.A(_03873_),
    .B(_01274_),
    .X(_03565_));
 sky130_fd_sc_hd__and2_1 _07428_ (.A(_03873_),
    .B(_01304_),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_1 _07429_ (.A(_03871_),
    .X(_03874_));
 sky130_fd_sc_hd__and2_1 _07430_ (.A(_03874_),
    .B(_01303_),
    .X(_03563_));
 sky130_fd_sc_hd__and2_1 _07431_ (.A(_03874_),
    .B(_01302_),
    .X(_03562_));
 sky130_fd_sc_hd__and2_1 _07432_ (.A(_03874_),
    .B(_01301_),
    .X(_03561_));
 sky130_fd_sc_hd__buf_1 _07433_ (.A(_03861_),
    .X(_03875_));
 sky130_fd_sc_hd__buf_1 _07434_ (.A(_03875_),
    .X(_03876_));
 sky130_fd_sc_hd__clkbuf_1 _07435_ (.A(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__and2_1 _07436_ (.A(_03877_),
    .B(_01300_),
    .X(_03560_));
 sky130_fd_sc_hd__and2_1 _07437_ (.A(_03877_),
    .B(_01299_),
    .X(_03559_));
 sky130_fd_sc_hd__and2_1 _07438_ (.A(_03877_),
    .B(_01298_),
    .X(_03558_));
 sky130_fd_sc_hd__clkbuf_1 _07439_ (.A(_03876_),
    .X(_03878_));
 sky130_fd_sc_hd__and2_1 _07440_ (.A(_03878_),
    .B(_01295_),
    .X(_03557_));
 sky130_fd_sc_hd__and2_1 _07441_ (.A(_03878_),
    .B(_01284_),
    .X(_03556_));
 sky130_fd_sc_hd__and2_1 _07442_ (.A(_03878_),
    .B(_01273_),
    .X(_03555_));
 sky130_fd_sc_hd__buf_1 _07443_ (.A(_03876_),
    .X(_03879_));
 sky130_fd_sc_hd__and2_1 _07444_ (.A(_03879_),
    .B(_01329_),
    .X(_03554_));
 sky130_fd_sc_hd__and2_1 _07445_ (.A(_03879_),
    .B(_01328_),
    .X(_03553_));
 sky130_fd_sc_hd__and2_1 _07446_ (.A(_03879_),
    .B(_01326_),
    .X(_03552_));
 sky130_fd_sc_hd__clkbuf_2 _07447_ (.A(_03875_),
    .X(_03880_));
 sky130_fd_sc_hd__clkbuf_1 _07448_ (.A(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__and2_1 _07449_ (.A(_03881_),
    .B(_01325_),
    .X(_03551_));
 sky130_fd_sc_hd__and2_1 _07450_ (.A(_03881_),
    .B(_01324_),
    .X(_03550_));
 sky130_fd_sc_hd__and2_1 _07451_ (.A(_03881_),
    .B(_01323_),
    .X(_03549_));
 sky130_fd_sc_hd__clkbuf_1 _07452_ (.A(_03880_),
    .X(_03882_));
 sky130_fd_sc_hd__and2_1 _07453_ (.A(_03882_),
    .B(_01322_),
    .X(_03548_));
 sky130_fd_sc_hd__and2_1 _07454_ (.A(_03882_),
    .B(_01321_),
    .X(_03547_));
 sky130_fd_sc_hd__and2_1 _07455_ (.A(_03882_),
    .B(_01320_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _07456_ (.A(_03880_),
    .X(_03883_));
 sky130_fd_sc_hd__and2_1 _07457_ (.A(_03883_),
    .B(_01319_),
    .X(_03545_));
 sky130_fd_sc_hd__and2_1 _07458_ (.A(_03883_),
    .B(_01318_),
    .X(_03544_));
 sky130_fd_sc_hd__and2_1 _07459_ (.A(_03883_),
    .B(_01317_),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_2 _07460_ (.A(_03875_),
    .X(_03884_));
 sky130_fd_sc_hd__clkbuf_1 _07461_ (.A(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__and2_1 _07462_ (.A(_03885_),
    .B(_01315_),
    .X(_03542_));
 sky130_fd_sc_hd__and2_1 _07463_ (.A(_03885_),
    .B(_01314_),
    .X(_03541_));
 sky130_fd_sc_hd__and2_1 _07464_ (.A(_03885_),
    .B(_01313_),
    .X(_03540_));
 sky130_fd_sc_hd__buf_1 _07465_ (.A(_03884_),
    .X(_03886_));
 sky130_fd_sc_hd__and2_1 _07466_ (.A(_03886_),
    .B(_01312_),
    .X(_03539_));
 sky130_fd_sc_hd__and2_1 _07467_ (.A(_03886_),
    .B(_01311_),
    .X(_03538_));
 sky130_fd_sc_hd__and2_1 _07468_ (.A(_03886_),
    .B(_01310_),
    .X(_03537_));
 sky130_fd_sc_hd__clkbuf_1 _07469_ (.A(_03884_),
    .X(_03887_));
 sky130_fd_sc_hd__and2_1 _07470_ (.A(_03887_),
    .B(_01309_),
    .X(_03536_));
 sky130_fd_sc_hd__and2_1 _07471_ (.A(_03887_),
    .B(_01308_),
    .X(_03535_));
 sky130_fd_sc_hd__and2_1 _07472_ (.A(_03887_),
    .B(_01307_),
    .X(_03534_));
 sky130_fd_sc_hd__buf_1 _07473_ (.A(_03861_),
    .X(_03888_));
 sky130_fd_sc_hd__buf_1 _07474_ (.A(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__buf_1 _07475_ (.A(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__and2_1 _07476_ (.A(_03890_),
    .B(_01306_),
    .X(_03533_));
 sky130_fd_sc_hd__and2_1 _07477_ (.A(_03890_),
    .B(_01336_),
    .X(_03532_));
 sky130_fd_sc_hd__and2_1 _07478_ (.A(_03890_),
    .B(_01335_),
    .X(_03531_));
 sky130_fd_sc_hd__clkbuf_1 _07479_ (.A(_03889_),
    .X(_03891_));
 sky130_fd_sc_hd__and2_1 _07480_ (.A(_03891_),
    .B(_01334_),
    .X(_03530_));
 sky130_fd_sc_hd__and2_1 _07481_ (.A(_03891_),
    .B(_01333_),
    .X(_03529_));
 sky130_fd_sc_hd__and2_1 _07482_ (.A(_03891_),
    .B(_01332_),
    .X(_03528_));
 sky130_fd_sc_hd__clkbuf_1 _07483_ (.A(_03889_),
    .X(_03892_));
 sky130_fd_sc_hd__and2_1 _07484_ (.A(_03892_),
    .B(_01331_),
    .X(_03527_));
 sky130_fd_sc_hd__and2_1 _07485_ (.A(_03892_),
    .B(_01330_),
    .X(_03526_));
 sky130_fd_sc_hd__and2_1 _07486_ (.A(_03892_),
    .B(_01327_),
    .X(_03525_));
 sky130_fd_sc_hd__buf_1 _07487_ (.A(_03888_),
    .X(_03893_));
 sky130_fd_sc_hd__buf_1 _07488_ (.A(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__and2_1 _07489_ (.A(_03894_),
    .B(_01316_),
    .X(_03524_));
 sky130_fd_sc_hd__and2_1 _07490_ (.A(_03894_),
    .B(_01305_),
    .X(_03523_));
 sky130_fd_sc_hd__nor2_1 _07491_ (.A(_03855_),
    .B(_03811_),
    .Y(_03521_));
 sky130_fd_sc_hd__buf_1 _07492_ (.A(_03854_),
    .X(_03895_));
 sky130_fd_sc_hd__nor2_1 _07493_ (.A(_03895_),
    .B(_03819_),
    .Y(_03520_));
 sky130_fd_sc_hd__nor2_1 _07494_ (.A(_03895_),
    .B(_03821_),
    .Y(_03519_));
 sky130_fd_sc_hd__nor2_1 _07495_ (.A(_03895_),
    .B(_03825_),
    .Y(_03518_));
 sky130_fd_sc_hd__buf_1 _07496_ (.A(_03854_),
    .X(_03896_));
 sky130_fd_sc_hd__nor2_1 _07497_ (.A(_03896_),
    .B(_03829_),
    .Y(_03517_));
 sky130_fd_sc_hd__nor2_1 _07498_ (.A(_03896_),
    .B(_03831_),
    .Y(_03516_));
 sky130_fd_sc_hd__inv_2 _07499_ (.A(\c1.instruction1[14] ),
    .Y(_03897_));
 sky130_fd_sc_hd__nor2_1 _07500_ (.A(_03896_),
    .B(_03897_),
    .Y(_03515_));
 sky130_fd_sc_hd__buf_1 _07501_ (.A(_03804_),
    .X(_03898_));
 sky130_fd_sc_hd__buf_1 _07502_ (.A(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__inv_2 _07503_ (.A(\c1.instruction1[13] ),
    .Y(_03900_));
 sky130_fd_sc_hd__nor2_1 _07504_ (.A(_03899_),
    .B(_03900_),
    .Y(_03514_));
 sky130_fd_sc_hd__nor2_1 _07505_ (.A(_03899_),
    .B(_03793_),
    .Y(_03513_));
 sky130_fd_sc_hd__nor2_1 _07506_ (.A(_03899_),
    .B(_03834_),
    .Y(_03512_));
 sky130_fd_sc_hd__buf_1 _07507_ (.A(_03898_),
    .X(_03901_));
 sky130_fd_sc_hd__nor2_1 _07508_ (.A(_03901_),
    .B(_03841_),
    .Y(_03511_));
 sky130_fd_sc_hd__nor2_1 _07509_ (.A(_03901_),
    .B(_03845_),
    .Y(_03510_));
 sky130_fd_sc_hd__nor2_1 _07510_ (.A(_03901_),
    .B(_03850_),
    .Y(_03509_));
 sky130_fd_sc_hd__buf_1 _07511_ (.A(_03898_),
    .X(_03902_));
 sky130_fd_sc_hd__nor2_1 _07512_ (.A(_03902_),
    .B(_03806_),
    .Y(_03508_));
 sky130_fd_sc_hd__nor2_1 _07513_ (.A(_03902_),
    .B(_03807_),
    .Y(_03507_));
 sky130_fd_sc_hd__nor2_1 _07514_ (.A(_03902_),
    .B(_03797_),
    .Y(_03506_));
 sky130_fd_sc_hd__clkbuf_1 _07515_ (.A(_03805_),
    .X(_03903_));
 sky130_fd_sc_hd__or2_1 _07516_ (.A(_03903_),
    .B(\c1.instruction1[4] ),
    .X(_03505_));
 sky130_fd_sc_hd__and2_1 _07517_ (.A(_03894_),
    .B(\c1.instruction1[3] ),
    .X(_03504_));
 sky130_fd_sc_hd__buf_1 _07518_ (.A(_03893_),
    .X(_03904_));
 sky130_fd_sc_hd__and2_1 _07519_ (.A(_03904_),
    .B(\c1.instruction1[2] ),
    .X(_03503_));
 sky130_fd_sc_hd__or2_1 _07520_ (.A(_03903_),
    .B(\c1.instruction1[1] ),
    .X(_03502_));
 sky130_fd_sc_hd__clkbuf_1 _07521_ (.A(_03805_),
    .X(_03905_));
 sky130_fd_sc_hd__or2_1 _07522_ (.A(_03905_),
    .B(\c1.instruction1[0] ),
    .X(_03501_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_opt_2_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__buf_1 _07524_ (.A(net56),
    .X(_03907_));
 sky130_fd_sc_hd__buf_1 _07525_ (.A(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__buf_1 _07526_ (.A(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__clkbuf_2 _07527_ (.A(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__buf_1 _07528_ (.A(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__clkbuf_2 _07529_ (.A(_03911_),
    .X(_02396_));
 sky130_fd_sc_hd__inv_2 _07530_ (.A(\c1.instruction3[11] ),
    .Y(_03912_));
 sky130_fd_sc_hd__inv_2 _07531_ (.A(\c1.instruction3[7] ),
    .Y(_03913_));
 sky130_fd_sc_hd__o22a_1 _07532_ (.A1(_03912_),
    .A2(net54),
    .B1(_03913_),
    .B2(net28),
    .X(_03914_));
 sky130_fd_sc_hd__inv_2 _07533_ (.A(net15),
    .Y(_03915_));
 sky130_fd_sc_hd__inv_2 _07534_ (.A(net54),
    .Y(_03916_));
 sky130_fd_sc_hd__inv_2 _07535_ (.A(\c1.instruction3[8] ),
    .Y(_03917_));
 sky130_fd_sc_hd__inv_2 _07536_ (.A(\c1.instruction1[18] ),
    .Y(_03918_));
 sky130_fd_sc_hd__o22a_1 _07537_ (.A1(_03917_),
    .A2(net20),
    .B1(\c1.instruction3[10] ),
    .B2(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__o221a_1 _07538_ (.A1(\c1.instruction3[9] ),
    .A2(_03915_),
    .B1(\c1.instruction3[11] ),
    .B2(_03916_),
    .C1(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__inv_2 _07539_ (.A(\c1.instruction3[9] ),
    .Y(_03921_));
 sky130_fd_sc_hd__inv_2 _07540_ (.A(\c1.instruction3[10] ),
    .Y(_03922_));
 sky130_fd_sc_hd__inv_2 _07541_ (.A(net20),
    .Y(_03923_));
 sky130_fd_sc_hd__inv_2 _07542_ (.A(net28),
    .Y(_03924_));
 sky130_fd_sc_hd__o22a_1 _07543_ (.A1(\c1.instruction3[8] ),
    .A2(_03923_),
    .B1(\c1.instruction3[7] ),
    .B2(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__o221a_1 _07544_ (.A1(_03921_),
    .A2(net15),
    .B1(_03922_),
    .B2(\c1.instruction1[18] ),
    .C1(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__and3_1 _07545_ (.A(_03914_),
    .B(_03920_),
    .C(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__inv_2 _07546_ (.A(\c1.instruction2[11] ),
    .Y(_03928_));
 sky130_fd_sc_hd__inv_2 _07547_ (.A(\c1.instruction2[7] ),
    .Y(_03929_));
 sky130_fd_sc_hd__o22a_1 _07548_ (.A1(_03928_),
    .A2(net54),
    .B1(_03929_),
    .B2(net28),
    .X(_03930_));
 sky130_fd_sc_hd__inv_2 _07549_ (.A(\c1.instruction2[8] ),
    .Y(_03931_));
 sky130_fd_sc_hd__o22a_1 _07550_ (.A1(_03931_),
    .A2(net20),
    .B1(\c1.instruction2[10] ),
    .B2(_03918_),
    .X(_03932_));
 sky130_fd_sc_hd__o221a_1 _07551_ (.A1(\c1.instruction2[9] ),
    .A2(_03915_),
    .B1(\c1.instruction2[11] ),
    .B2(_03916_),
    .C1(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__inv_2 _07552_ (.A(\c1.instruction2[9] ),
    .Y(_03934_));
 sky130_fd_sc_hd__inv_2 _07553_ (.A(\c1.instruction2[10] ),
    .Y(_03935_));
 sky130_fd_sc_hd__o22a_1 _07554_ (.A1(\c1.instruction2[8] ),
    .A2(_03923_),
    .B1(\c1.instruction2[7] ),
    .B2(_03924_),
    .X(_03936_));
 sky130_fd_sc_hd__o221a_1 _07555_ (.A1(_03934_),
    .A2(net15),
    .B1(_03935_),
    .B2(\c1.instruction1[18] ),
    .C1(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__and3_1 _07556_ (.A(_03930_),
    .B(_03933_),
    .C(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__o21ba_1 _07557_ (.A1(_03927_),
    .A2(_03938_),
    .B1_N(_03790_),
    .X(_03939_));
 sky130_fd_sc_hd__inv_2 _07558_ (.A(_03927_),
    .Y(_03940_));
 sky130_fd_sc_hd__or4_4 _07559_ (.A(_03788_),
    .B(_03789_),
    .C(_03787_),
    .D(_03797_),
    .X(_03941_));
 sky130_fd_sc_hd__o211ai_2 _07560_ (.A1(_03801_),
    .A2(_03940_),
    .B1(_03823_),
    .C1(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__o22a_1 _07561_ (.A1(net50),
    .A2(_03913_),
    .B1(_03842_),
    .B2(\c1.instruction3[10] ),
    .X(_03943_));
 sky130_fd_sc_hd__o221a_1 _07562_ (.A1(_03857_),
    .A2(\c1.instruction3[7] ),
    .B1(\c1.instruction1[22] ),
    .B2(_03921_),
    .C1(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__o22a_1 _07563_ (.A1(_03836_),
    .A2(\c1.instruction3[11] ),
    .B1(_03851_),
    .B2(\c1.instruction3[8] ),
    .X(_03945_));
 sky130_fd_sc_hd__o221a_1 _07564_ (.A1(net53),
    .A2(_03912_),
    .B1(\c1.instruction1[23] ),
    .B2(_03922_),
    .C1(_03945_),
    .X(_03946_));
 sky130_fd_sc_hd__o221a_1 _07565_ (.A1(net40),
    .A2(_03917_),
    .B1(_03846_),
    .B2(\c1.instruction3[9] ),
    .C1(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__o211a_1 _07566_ (.A1(_03939_),
    .A2(_03942_),
    .B1(_03944_),
    .C1(_03947_),
    .X(_03500_));
 sky130_fd_sc_hd__and2_1 _07567_ (.A(_03904_),
    .B(\e1.alu1.out[31] ),
    .X(_03499_));
 sky130_fd_sc_hd__and2_1 _07568_ (.A(_03904_),
    .B(\e1.alu1.out[30] ),
    .X(_03498_));
 sky130_fd_sc_hd__clkbuf_2 _07569_ (.A(_03893_),
    .X(_03948_));
 sky130_fd_sc_hd__and2_1 _07570_ (.A(_03948_),
    .B(\e1.alu1.out[29] ),
    .X(_03497_));
 sky130_fd_sc_hd__and2_1 _07571_ (.A(_03948_),
    .B(\e1.alu1.out[28] ),
    .X(_03496_));
 sky130_fd_sc_hd__and2_1 _07572_ (.A(_03948_),
    .B(\e1.alu1.out[27] ),
    .X(_03495_));
 sky130_fd_sc_hd__clkbuf_2 _07573_ (.A(_03888_),
    .X(_03949_));
 sky130_fd_sc_hd__buf_1 _07574_ (.A(_03949_),
    .X(_03950_));
 sky130_fd_sc_hd__and2_1 _07575_ (.A(_03950_),
    .B(\e1.alu1.out[26] ),
    .X(_03494_));
 sky130_fd_sc_hd__and2_1 _07576_ (.A(_03950_),
    .B(\e1.alu1.out[25] ),
    .X(_03493_));
 sky130_fd_sc_hd__and2_1 _07577_ (.A(_03950_),
    .B(\e1.alu1.out[24] ),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_1 _07578_ (.A(_03949_),
    .X(_03951_));
 sky130_fd_sc_hd__and2_1 _07579_ (.A(_03951_),
    .B(\e1.alu1.out[23] ),
    .X(_03491_));
 sky130_fd_sc_hd__and2_1 _07580_ (.A(_03951_),
    .B(\e1.alu1.out[22] ),
    .X(_03490_));
 sky130_fd_sc_hd__and2_1 _07581_ (.A(_03951_),
    .B(\e1.alu1.out[21] ),
    .X(_03489_));
 sky130_fd_sc_hd__clkbuf_1 _07582_ (.A(_03949_),
    .X(_03952_));
 sky130_fd_sc_hd__and2_1 _07583_ (.A(_03952_),
    .B(\e1.alu1.out[20] ),
    .X(_03488_));
 sky130_fd_sc_hd__and2_1 _07584_ (.A(_03952_),
    .B(\e1.alu1.out[19] ),
    .X(_03487_));
 sky130_fd_sc_hd__and2_1 _07585_ (.A(_03952_),
    .B(\e1.alu1.out[18] ),
    .X(_03486_));
 sky130_fd_sc_hd__buf_1 _07586_ (.A(_03666_),
    .X(_03953_));
 sky130_fd_sc_hd__buf_1 _07587_ (.A(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__buf_1 _07588_ (.A(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__and2_1 _07589_ (.A(_03955_),
    .B(\e1.alu1.out[17] ),
    .X(_03485_));
 sky130_fd_sc_hd__and2_1 _07590_ (.A(_03955_),
    .B(\e1.alu1.out[16] ),
    .X(_03484_));
 sky130_fd_sc_hd__and2_1 _07591_ (.A(_03955_),
    .B(\e1.alu1.out[15] ),
    .X(_03483_));
 sky130_fd_sc_hd__clkbuf_1 _07592_ (.A(_03954_),
    .X(_03956_));
 sky130_fd_sc_hd__and2_1 _07593_ (.A(_03956_),
    .B(\e1.alu1.out[14] ),
    .X(_03482_));
 sky130_fd_sc_hd__and2_1 _07594_ (.A(_03956_),
    .B(\e1.alu1.out[13] ),
    .X(_03481_));
 sky130_fd_sc_hd__and2_1 _07595_ (.A(_03956_),
    .B(\e1.alu1.out[12] ),
    .X(_03480_));
 sky130_fd_sc_hd__buf_1 _07596_ (.A(_03954_),
    .X(_03957_));
 sky130_fd_sc_hd__and2_1 _07597_ (.A(_03957_),
    .B(\e1.alu1.out[11] ),
    .X(_03479_));
 sky130_fd_sc_hd__and2_1 _07598_ (.A(_03957_),
    .B(\e1.alu1.out[10] ),
    .X(_03478_));
 sky130_fd_sc_hd__and2_1 _07599_ (.A(_03957_),
    .B(\e1.alu1.out[9] ),
    .X(_03477_));
 sky130_fd_sc_hd__buf_1 _07600_ (.A(_03953_),
    .X(_03958_));
 sky130_fd_sc_hd__clkbuf_1 _07601_ (.A(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__and2_1 _07602_ (.A(_03959_),
    .B(\e1.alu1.out[8] ),
    .X(_03476_));
 sky130_fd_sc_hd__and2_1 _07603_ (.A(_03959_),
    .B(\e1.alu1.out[7] ),
    .X(_03475_));
 sky130_fd_sc_hd__and2_1 _07604_ (.A(_03959_),
    .B(\e1.alu1.out[6] ),
    .X(_03474_));
 sky130_fd_sc_hd__clkbuf_1 _07605_ (.A(_03958_),
    .X(_03960_));
 sky130_fd_sc_hd__and2_1 _07606_ (.A(_03960_),
    .B(\e1.alu1.out[5] ),
    .X(_03473_));
 sky130_fd_sc_hd__and2_1 _07607_ (.A(_03960_),
    .B(\e1.alu1.out[4] ),
    .X(_03472_));
 sky130_fd_sc_hd__and2_1 _07608_ (.A(_03960_),
    .B(\e1.alu1.out[3] ),
    .X(_03471_));
 sky130_fd_sc_hd__buf_1 _07609_ (.A(_03958_),
    .X(_03961_));
 sky130_fd_sc_hd__and2_1 _07610_ (.A(_03961_),
    .B(\e1.alu1.out[2] ),
    .X(_03470_));
 sky130_fd_sc_hd__and2_1 _07611_ (.A(_03961_),
    .B(\e1.alu1.out[1] ),
    .X(_03469_));
 sky130_fd_sc_hd__and2_1 _07612_ (.A(_03864_),
    .B(\e1.alu1.out[0] ),
    .X(_03468_));
 sky130_fd_sc_hd__buf_1 _07613_ (.A(_03804_),
    .X(_03962_));
 sky130_fd_sc_hd__buf_1 _07614_ (.A(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__buf_1 _07615_ (.A(\c1.instruction2[14] ),
    .X(_03964_));
 sky130_fd_sc_hd__inv_2 _07616_ (.A(_03964_),
    .Y(_03965_));
 sky130_fd_sc_hd__buf_1 _07617_ (.A(_03965_),
    .X(_03966_));
 sky130_fd_sc_hd__buf_1 _07618_ (.A(_03966_),
    .X(_00004_));
 sky130_fd_sc_hd__nor2_1 _07619_ (.A(_03963_),
    .B(_00004_),
    .Y(_03467_));
 sky130_fd_sc_hd__inv_2 _07620_ (.A(\c1.instruction2[13] ),
    .Y(_03967_));
 sky130_fd_sc_hd__buf_1 _07621_ (.A(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__buf_1 _07622_ (.A(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__nor2_1 _07623_ (.A(_03963_),
    .B(_03969_),
    .Y(_03466_));
 sky130_fd_sc_hd__inv_2 _07624_ (.A(\c1.instruction2[12] ),
    .Y(_03970_));
 sky130_fd_sc_hd__buf_1 _07625_ (.A(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__nor2_1 _07626_ (.A(_03963_),
    .B(_03971_),
    .Y(_03465_));
 sky130_fd_sc_hd__buf_1 _07627_ (.A(_03962_),
    .X(_03972_));
 sky130_fd_sc_hd__nor2_1 _07628_ (.A(_03972_),
    .B(_03928_),
    .Y(_03464_));
 sky130_fd_sc_hd__nor2_1 _07629_ (.A(_03972_),
    .B(_03935_),
    .Y(_03463_));
 sky130_fd_sc_hd__nor2_1 _07630_ (.A(_03972_),
    .B(_03934_),
    .Y(_03462_));
 sky130_fd_sc_hd__buf_1 _07631_ (.A(_03962_),
    .X(_03973_));
 sky130_fd_sc_hd__nor2_1 _07632_ (.A(_03973_),
    .B(_03931_),
    .Y(_03461_));
 sky130_fd_sc_hd__nor2_1 _07633_ (.A(_03973_),
    .B(_03929_),
    .Y(_03460_));
 sky130_fd_sc_hd__nor2_1 _07634_ (.A(_03973_),
    .B(_03676_),
    .Y(_03459_));
 sky130_fd_sc_hd__nor2_1 _07635_ (.A(_03903_),
    .B(_03677_),
    .Y(_03458_));
 sky130_fd_sc_hd__buf_1 _07636_ (.A(\c1.instruction2[4] ),
    .X(_03974_));
 sky130_fd_sc_hd__or2_1 _07637_ (.A(_03905_),
    .B(_03974_),
    .X(_03457_));
 sky130_fd_sc_hd__and2_1 _07638_ (.A(_03961_),
    .B(\c1.instruction2[3] ),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_2 _07639_ (.A(_03673_),
    .X(_03975_));
 sky130_fd_sc_hd__and2_1 _07640_ (.A(_03975_),
    .B(\c1.instruction2[2] ),
    .X(_03455_));
 sky130_fd_sc_hd__or2_1 _07641_ (.A(_03905_),
    .B(\c1.instruction2[1] ),
    .X(_03454_));
 sky130_fd_sc_hd__or2_1 _07642_ (.A(_03665_),
    .B(\c1.instruction2[0] ),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_2 _07643_ (.A(\e1.offset[11] ),
    .X(_03976_));
 sky130_fd_sc_hd__inv_2 _07644_ (.A(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__buf_1 _07645_ (.A(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__clkbuf_1 _07646_ (.A(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__buf_1 _07647_ (.A(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__buf_1 _07648_ (.A(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__clkbuf_1 _07649_ (.A(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__buf_1 _07650_ (.A(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__clkbuf_1 _07651_ (.A(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__buf_1 _07652_ (.A(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__buf_1 _07653_ (.A(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__clkbuf_1 _07654_ (.A(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__buf_1 _07655_ (.A(_03987_),
    .X(_03988_));
 sky130_fd_sc_hd__buf_1 _07656_ (.A(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__buf_1 _07657_ (.A(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__buf_1 _07658_ (.A(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__buf_1 _07659_ (.A(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__buf_1 _07660_ (.A(_03976_),
    .X(_03993_));
 sky130_fd_sc_hd__inv_2 _07661_ (.A(_01271_),
    .Y(_03994_));
 sky130_fd_sc_hd__o22a_1 _07662_ (.A1(_03990_),
    .A2(_01271_),
    .B1(_03993_),
    .B2(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__clkbuf_1 _07663_ (.A(_03988_),
    .X(_03996_));
 sky130_fd_sc_hd__buf_1 _07664_ (.A(_01267_),
    .X(_03997_));
 sky130_fd_sc_hd__a2bb2o_1 _07665_ (.A1_N(_03996_),
    .A2_N(_03997_),
    .B1(_03996_),
    .B2(_01267_),
    .X(_03998_));
 sky130_fd_sc_hd__inv_2 _07666_ (.A(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__a2bb2o_1 _07667_ (.A1_N(_03996_),
    .A2_N(_01269_),
    .B1(_03988_),
    .B2(_01269_),
    .X(_04000_));
 sky130_fd_sc_hd__inv_2 _07668_ (.A(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__clkbuf_1 _07669_ (.A(_03986_),
    .X(_04002_));
 sky130_fd_sc_hd__clkbuf_1 _07670_ (.A(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__buf_1 _07671_ (.A(_01263_),
    .X(_04004_));
 sky130_fd_sc_hd__a2bb2o_1 _07672_ (.A1_N(_04003_),
    .A2_N(_04004_),
    .B1(_04003_),
    .B2(_01263_),
    .X(_04005_));
 sky130_fd_sc_hd__a2bb2o_1 _07673_ (.A1_N(_03987_),
    .A2_N(_01265_),
    .B1(_03987_),
    .B2(_01265_),
    .X(_04006_));
 sky130_fd_sc_hd__buf_1 _07674_ (.A(_01259_),
    .X(_04007_));
 sky130_fd_sc_hd__clkbuf_1 _07675_ (.A(_03986_),
    .X(_04008_));
 sky130_fd_sc_hd__a2bb2o_1 _07676_ (.A1_N(_04002_),
    .A2_N(_04007_),
    .B1(_04008_),
    .B2(_01259_),
    .X(_04009_));
 sky130_fd_sc_hd__a2bb2o_1 _07677_ (.A1_N(_04008_),
    .A2_N(_01261_),
    .B1(_04008_),
    .B2(_01261_),
    .X(_04010_));
 sky130_fd_sc_hd__buf_1 _07678_ (.A(_01243_),
    .X(_04011_));
 sky130_fd_sc_hd__clkbuf_1 _07679_ (.A(_03978_),
    .X(_04012_));
 sky130_fd_sc_hd__buf_1 _07680_ (.A(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__or2_1 _07681_ (.A(_04013_),
    .B(_01245_),
    .X(_04014_));
 sky130_fd_sc_hd__buf_1 _07682_ (.A(_03983_),
    .X(_04015_));
 sky130_fd_sc_hd__buf_1 _07683_ (.A(_01247_),
    .X(_04016_));
 sky130_fd_sc_hd__o22a_1 _07684_ (.A1(_04015_),
    .A2(_04016_),
    .B1(_04015_),
    .B2(_01249_),
    .X(_04017_));
 sky130_fd_sc_hd__o211a_1 _07685_ (.A1(_03985_),
    .A2(_04011_),
    .B1(_04014_),
    .C1(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__buf_1 _07686_ (.A(_01253_),
    .X(_04019_));
 sky130_fd_sc_hd__or2_2 _07687_ (.A(_03980_),
    .B(_01251_),
    .X(_04020_));
 sky130_fd_sc_hd__buf_1 _07688_ (.A(_01255_),
    .X(_04021_));
 sky130_fd_sc_hd__clkbuf_1 _07689_ (.A(_03983_),
    .X(_04022_));
 sky130_fd_sc_hd__o22a_1 _07690_ (.A1(_04015_),
    .A2(_04021_),
    .B1(_04022_),
    .B2(_01257_),
    .X(_04023_));
 sky130_fd_sc_hd__o211a_1 _07691_ (.A1(_03985_),
    .A2(_04019_),
    .B1(_04020_),
    .C1(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__a2bb2o_1 _07692_ (.A1_N(_04022_),
    .A2_N(_04021_),
    .B1(_04022_),
    .B2(_01255_),
    .X(_04025_));
 sky130_fd_sc_hd__a2bb2o_1 _07693_ (.A1_N(_03984_),
    .A2_N(_01257_),
    .B1(_03984_),
    .B2(_01257_),
    .X(_04026_));
 sky130_fd_sc_hd__buf_1 _07694_ (.A(_03981_),
    .X(_04027_));
 sky130_fd_sc_hd__inv_2 _07695_ (.A(_04020_),
    .Y(_04028_));
 sky130_fd_sc_hd__a21oi_2 _07696_ (.A1(_04027_),
    .A2(_01251_),
    .B1(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__inv_2 _07697_ (.A(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__a2bb2o_1 _07698_ (.A1_N(_04027_),
    .A2_N(_04019_),
    .B1(_04027_),
    .B2(_01253_),
    .X(_04031_));
 sky130_fd_sc_hd__or2_1 _07699_ (.A(_04030_),
    .B(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__a2bb2o_1 _07700_ (.A1_N(_03982_),
    .A2_N(_01243_),
    .B1(_03982_),
    .B2(_01243_),
    .X(_04033_));
 sky130_fd_sc_hd__clkbuf_1 _07701_ (.A(_03981_),
    .X(_04034_));
 sky130_fd_sc_hd__a21bo_1 _07702_ (.A1(_04034_),
    .A2(_01245_),
    .B1_N(_04014_),
    .X(_04035_));
 sky130_fd_sc_hd__or2_1 _07703_ (.A(_04033_),
    .B(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__a2bb2o_1 _07704_ (.A1_N(_04034_),
    .A2_N(_01249_),
    .B1(_04034_),
    .B2(_01249_),
    .X(_04037_));
 sky130_fd_sc_hd__inv_2 _07705_ (.A(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__buf_1 _07706_ (.A(_04013_),
    .X(_04039_));
 sky130_fd_sc_hd__a2bb2o_1 _07707_ (.A1_N(_04039_),
    .A2_N(_04016_),
    .B1(_04039_),
    .B2(_01247_),
    .X(_04040_));
 sky130_fd_sc_hd__inv_2 _07708_ (.A(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__buf_1 _07709_ (.A(_01235_),
    .X(_04042_));
 sky130_fd_sc_hd__or2_1 _07710_ (.A(_03977_),
    .B(_01237_),
    .X(_04043_));
 sky130_fd_sc_hd__buf_1 _07711_ (.A(_01239_),
    .X(_04044_));
 sky130_fd_sc_hd__o22a_1 _07712_ (.A1(_04013_),
    .A2(_04044_),
    .B1(_03980_),
    .B2(_01241_),
    .X(_04045_));
 sky130_fd_sc_hd__a2bb2o_1 _07713_ (.A1_N(_04012_),
    .A2_N(_04044_),
    .B1(_04012_),
    .B2(_01239_),
    .X(_04046_));
 sky130_fd_sc_hd__a2bb2o_1 _07714_ (.A1_N(_03979_),
    .A2_N(_01241_),
    .B1(_03979_),
    .B2(_01241_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_1 _07715_ (.A(_03977_),
    .X(_04048_));
 sky130_fd_sc_hd__a2bb2o_1 _07716_ (.A1_N(_04048_),
    .A2_N(_01235_),
    .B1(_04048_),
    .B2(_01235_),
    .X(_04049_));
 sky130_fd_sc_hd__a21bo_1 _07717_ (.A1(_04048_),
    .A2(_01237_),
    .B1_N(_04043_),
    .X(_04050_));
 sky130_fd_sc_hd__or2_1 _07718_ (.A(_04049_),
    .B(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__inv_2 _07719_ (.A(_01233_),
    .Y(_04052_));
 sky130_fd_sc_hd__nor2_1 _07720_ (.A(_04052_),
    .B(\e1.offset[11] ),
    .Y(_04053_));
 sky130_fd_sc_hd__a21oi_2 _07721_ (.A1(_04052_),
    .A2(_03976_),
    .B1(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__inv_2 _07722_ (.A(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__buf_1 _07723_ (.A(_01231_),
    .X(_04056_));
 sky130_fd_sc_hd__inv_2 _07724_ (.A(\e1.offset[10] ),
    .Y(_04057_));
 sky130_fd_sc_hd__buf_1 _07725_ (.A(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__a2bb2o_1 _07726_ (.A1_N(_04056_),
    .A2_N(_04058_),
    .B1(_01231_),
    .B2(_04057_),
    .X(_04059_));
 sky130_fd_sc_hd__inv_2 _07727_ (.A(\e1.offset[9] ),
    .Y(_04060_));
 sky130_fd_sc_hd__nor2_1 _07728_ (.A(_01229_),
    .B(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__inv_2 _07729_ (.A(\e1.offset[8] ),
    .Y(_04062_));
 sky130_fd_sc_hd__nor2_1 _07730_ (.A(_01227_),
    .B(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__buf_1 _07731_ (.A(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__o2bb2a_1 _07732_ (.A1_N(_01229_),
    .A2_N(_04060_),
    .B1(_04061_),
    .B2(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__inv_2 _07733_ (.A(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__o32a_1 _07734_ (.A1(_04056_),
    .A2(_04058_),
    .A3(_04053_),
    .B1(_01233_),
    .B2(_03978_),
    .X(_04067_));
 sky130_fd_sc_hd__a21oi_1 _07735_ (.A1(_01229_),
    .A2(_04060_),
    .B1(_04061_),
    .Y(_04068_));
 sky130_fd_sc_hd__a21oi_1 _07736_ (.A1(_01227_),
    .A2(_04062_),
    .B1(_04063_),
    .Y(_04069_));
 sky130_fd_sc_hd__nand2_1 _07737_ (.A(_04068_),
    .B(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__inv_2 _07738_ (.A(_01225_),
    .Y(_04071_));
 sky130_fd_sc_hd__clkbuf_1 _07739_ (.A(_04071_),
    .X(_04072_));
 sky130_fd_sc_hd__clkbuf_1 _07740_ (.A(\e1.offset[7] ),
    .X(_04073_));
 sky130_fd_sc_hd__o2bb2a_1 _07741_ (.A1_N(_04072_),
    .A2_N(_04073_),
    .B1(_04072_),
    .B2(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__inv_2 _07742_ (.A(\e1.offset[6] ),
    .Y(_04075_));
 sky130_fd_sc_hd__inv_2 _07743_ (.A(_01223_),
    .Y(_04076_));
 sky130_fd_sc_hd__o22a_1 _07744_ (.A1(_01223_),
    .A2(_04075_),
    .B1(_04076_),
    .B2(\e1.offset[6] ),
    .X(_04077_));
 sky130_fd_sc_hd__inv_2 _07745_ (.A(_01221_),
    .Y(_04078_));
 sky130_fd_sc_hd__nor2_1 _07746_ (.A(_04078_),
    .B(\e1.offset[5] ),
    .Y(_04079_));
 sky130_fd_sc_hd__a21oi_2 _07747_ (.A1(_04078_),
    .A2(\e1.offset[5] ),
    .B1(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__clkbuf_1 _07748_ (.A(_01219_),
    .X(_04081_));
 sky130_fd_sc_hd__inv_2 _07749_ (.A(\e1.offset[4] ),
    .Y(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _07750_ (.A(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__a2bb2o_1 _07751_ (.A1_N(_04081_),
    .A2_N(_04083_),
    .B1(_04081_),
    .B2(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__inv_2 _07752_ (.A(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__inv_2 _07753_ (.A(_01217_),
    .Y(_04086_));
 sky130_fd_sc_hd__nor2_1 _07754_ (.A(_04086_),
    .B(\e1.offset[3] ),
    .Y(_04087_));
 sky130_fd_sc_hd__inv_2 _07755_ (.A(_01215_),
    .Y(_04088_));
 sky130_fd_sc_hd__nor2_1 _07756_ (.A(_04088_),
    .B(\e1.offset[2] ),
    .Y(_04089_));
 sky130_fd_sc_hd__inv_2 _07757_ (.A(\e1.offset[1] ),
    .Y(_04090_));
 sky130_fd_sc_hd__inv_2 _07758_ (.A(\e1.offset[0] ),
    .Y(_04091_));
 sky130_fd_sc_hd__a2bb2o_1 _07759_ (.A1_N(_01213_),
    .A2_N(_04090_),
    .B1(_01213_),
    .B2(_04090_),
    .X(_04092_));
 sky130_fd_sc_hd__or3_1 _07760_ (.A(_01211_),
    .B(_04091_),
    .C(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__o21ai_2 _07761_ (.A1(_01213_),
    .A2(_04090_),
    .B1(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__inv_2 _07762_ (.A(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__o2bb2a_1 _07763_ (.A1_N(_04088_),
    .A2_N(\e1.offset[2] ),
    .B1(_04089_),
    .B2(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__o2bb2a_1 _07764_ (.A1_N(_04086_),
    .A2_N(\e1.offset[3] ),
    .B1(_04087_),
    .B2(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__inv_2 _07765_ (.A(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__or3_2 _07766_ (.A(_01219_),
    .B(_04082_),
    .C(_04079_),
    .X(_04099_));
 sky130_fd_sc_hd__a21bo_1 _07767_ (.A1(_04078_),
    .A2(\e1.offset[5] ),
    .B1_N(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__a31o_1 _07768_ (.A1(_04080_),
    .A2(_04085_),
    .A3(_04098_),
    .B1(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__or2_1 _07769_ (.A(_04071_),
    .B(\e1.offset[7] ),
    .X(_04102_));
 sky130_fd_sc_hd__a32o_1 _07770_ (.A1(_04076_),
    .A2(\e1.offset[6] ),
    .A3(_04102_),
    .B1(_04072_),
    .B2(_04073_),
    .X(_04103_));
 sky130_fd_sc_hd__a31o_1 _07771_ (.A1(_04074_),
    .A2(_04077_),
    .A3(_04101_),
    .B1(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__or4b_4 _07772_ (.A(_04055_),
    .B(_04059_),
    .C(_04070_),
    .D_N(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__o311a_1 _07773_ (.A1(_04055_),
    .A2(_04059_),
    .A3(_04066_),
    .B1(_04067_),
    .C1(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__or4_4 _07774_ (.A(_04046_),
    .B(_04047_),
    .C(_04051_),
    .D(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__o2111a_1 _07775_ (.A1(_04039_),
    .A2(_04042_),
    .B1(_04043_),
    .C1(_04045_),
    .D1(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__inv_2 _07776_ (.A(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__and4b_1 _07777_ (.A_N(_04036_),
    .B(_04038_),
    .C(_04041_),
    .D(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__or4b_1 _07778_ (.A(_04025_),
    .B(_04026_),
    .C(_04032_),
    .D_N(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__and3_1 _07779_ (.A(_04018_),
    .B(_04024_),
    .C(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__or3_1 _07780_ (.A(_04009_),
    .B(_04010_),
    .C(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__buf_1 _07781_ (.A(_04002_),
    .X(_04114_));
 sky130_fd_sc_hd__o22a_1 _07782_ (.A1(_04114_),
    .A2(_04007_),
    .B1(_04003_),
    .B2(_01261_),
    .X(_04115_));
 sky130_fd_sc_hd__o22a_1 _07783_ (.A1(_04114_),
    .A2(_04004_),
    .B1(_04114_),
    .B2(_01265_),
    .X(_04116_));
 sky130_fd_sc_hd__o311a_1 _07784_ (.A1(_04005_),
    .A2(_04006_),
    .A3(_04113_),
    .B1(_04115_),
    .C1(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__inv_2 _07785_ (.A(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__buf_1 _07786_ (.A(_03989_),
    .X(_04119_));
 sky130_fd_sc_hd__o22ai_1 _07787_ (.A1(_03990_),
    .A2(_03997_),
    .B1(_04119_),
    .B2(_01269_),
    .Y(_04120_));
 sky130_fd_sc_hd__a31o_1 _07788_ (.A1(_03999_),
    .A2(_04001_),
    .A3(_04118_),
    .B1(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__nand2_1 _07789_ (.A(_03995_),
    .B(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__o21ai_1 _07790_ (.A1(_03992_),
    .A2(_01271_),
    .B1(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__a2bb2o_1 _07791_ (.A1_N(_03993_),
    .A2_N(_01272_),
    .B1(_03993_),
    .B2(_01272_),
    .X(_04124_));
 sky130_fd_sc_hd__inv_2 _07792_ (.A(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__inv_2 _07793_ (.A(_04123_),
    .Y(_04126_));
 sky130_fd_sc_hd__o221a_1 _07794_ (.A1(_04123_),
    .A2(_04125_),
    .B1(_04126_),
    .B2(_04124_),
    .C1(_03975_),
    .X(_03452_));
 sky130_fd_sc_hd__buf_1 _07795_ (.A(_03667_),
    .X(_04127_));
 sky130_fd_sc_hd__buf_1 _07796_ (.A(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__o211a_1 _07797_ (.A1(_03995_),
    .A2(_04121_),
    .B1(_04128_),
    .C1(_04122_),
    .X(_03451_));
 sky130_fd_sc_hd__or2_1 _07798_ (.A(_04117_),
    .B(_03998_),
    .X(_04129_));
 sky130_fd_sc_hd__o21ai_1 _07799_ (.A1(_03992_),
    .A2(_03997_),
    .B1(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__inv_2 _07800_ (.A(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__o221a_1 _07801_ (.A1(_04000_),
    .A2(_04131_),
    .B1(_04001_),
    .B2(_04130_),
    .C1(_03975_),
    .X(_03450_));
 sky130_fd_sc_hd__o211a_1 _07802_ (.A1(_04118_),
    .A2(_03999_),
    .B1(_04128_),
    .C1(_04129_),
    .X(_03449_));
 sky130_fd_sc_hd__inv_2 _07803_ (.A(_04005_),
    .Y(_04132_));
 sky130_fd_sc_hd__nand2_1 _07804_ (.A(_04113_),
    .B(_04115_),
    .Y(_04133_));
 sky130_fd_sc_hd__nand2_1 _07805_ (.A(_04132_),
    .B(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__o21ai_1 _07806_ (.A1(_03992_),
    .A2(_04004_),
    .B1(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__inv_2 _07807_ (.A(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__inv_2 _07808_ (.A(_04006_),
    .Y(_04137_));
 sky130_fd_sc_hd__buf_1 _07809_ (.A(_03953_),
    .X(_04138_));
 sky130_fd_sc_hd__buf_1 _07810_ (.A(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__o221a_1 _07811_ (.A1(_04006_),
    .A2(_04136_),
    .B1(_04137_),
    .B2(_04135_),
    .C1(_04139_),
    .X(_03448_));
 sky130_fd_sc_hd__o211a_1 _07812_ (.A1(_04132_),
    .A2(_04133_),
    .B1(_04128_),
    .C1(_04134_),
    .X(_03447_));
 sky130_fd_sc_hd__buf_1 _07813_ (.A(_03991_),
    .X(_04140_));
 sky130_fd_sc_hd__or2_1 _07814_ (.A(_04112_),
    .B(_04009_),
    .X(_04141_));
 sky130_fd_sc_hd__o21ai_1 _07815_ (.A1(_04140_),
    .A2(_04007_),
    .B1(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__inv_2 _07816_ (.A(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__inv_2 _07817_ (.A(_04010_),
    .Y(_04144_));
 sky130_fd_sc_hd__o221a_1 _07818_ (.A1(_04010_),
    .A2(_04143_),
    .B1(_04144_),
    .B2(_04142_),
    .C1(_04139_),
    .X(_03446_));
 sky130_fd_sc_hd__nand2_1 _07819_ (.A(_04112_),
    .B(_04009_),
    .Y(_04145_));
 sky130_fd_sc_hd__and3_1 _07820_ (.A(_03674_),
    .B(_04141_),
    .C(_04145_),
    .X(_03445_));
 sky130_fd_sc_hd__or2b_1 _07821_ (.A(_04110_),
    .B_N(_04018_),
    .X(_04146_));
 sky130_fd_sc_hd__inv_2 _07822_ (.A(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__o221a_1 _07823_ (.A1(_04119_),
    .A2(_04019_),
    .B1(_04032_),
    .B2(_04147_),
    .C1(_04020_),
    .X(_04148_));
 sky130_fd_sc_hd__or2_1 _07824_ (.A(_04025_),
    .B(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__o21ai_1 _07825_ (.A1(_04140_),
    .A2(_04021_),
    .B1(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__inv_2 _07826_ (.A(_04150_),
    .Y(_04151_));
 sky130_fd_sc_hd__inv_2 _07827_ (.A(_04026_),
    .Y(_04152_));
 sky130_fd_sc_hd__o221a_1 _07828_ (.A1(_04026_),
    .A2(_04151_),
    .B1(_04152_),
    .B2(_04150_),
    .C1(_04139_),
    .X(_03444_));
 sky130_fd_sc_hd__buf_1 _07829_ (.A(_04127_),
    .X(_04153_));
 sky130_fd_sc_hd__nand2_1 _07830_ (.A(_04025_),
    .B(_04148_),
    .Y(_04154_));
 sky130_fd_sc_hd__and3_1 _07831_ (.A(_04153_),
    .B(_04149_),
    .C(_04154_),
    .X(_03443_));
 sky130_fd_sc_hd__or2_1 _07832_ (.A(_04030_),
    .B(_04147_),
    .X(_04155_));
 sky130_fd_sc_hd__inv_2 _07833_ (.A(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__inv_2 _07834_ (.A(_04031_),
    .Y(_04157_));
 sky130_fd_sc_hd__buf_1 _07835_ (.A(_03673_),
    .X(_04158_));
 sky130_fd_sc_hd__o21ai_1 _07836_ (.A1(_04028_),
    .A2(_04156_),
    .B1(_04157_),
    .Y(_04159_));
 sky130_fd_sc_hd__o311a_1 _07837_ (.A1(_04028_),
    .A2(_04156_),
    .A3(_04157_),
    .B1(_04158_),
    .C1(_04159_),
    .X(_03442_));
 sky130_fd_sc_hd__buf_1 _07838_ (.A(_04127_),
    .X(_04160_));
 sky130_fd_sc_hd__o211a_1 _07839_ (.A1(_04029_),
    .A2(_04146_),
    .B1(_04160_),
    .C1(_04155_),
    .X(_03441_));
 sky130_fd_sc_hd__o221a_1 _07840_ (.A1(_04119_),
    .A2(_04011_),
    .B1(_04108_),
    .B2(_04036_),
    .C1(_04014_),
    .X(_04161_));
 sky130_fd_sc_hd__or2_1 _07841_ (.A(_04040_),
    .B(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__o21ai_1 _07842_ (.A1(_04140_),
    .A2(_04016_),
    .B1(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__inv_2 _07843_ (.A(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__buf_1 _07844_ (.A(_04138_),
    .X(_04165_));
 sky130_fd_sc_hd__o221a_1 _07845_ (.A1(_04037_),
    .A2(_04164_),
    .B1(_04038_),
    .B2(_04163_),
    .C1(_04165_),
    .X(_03440_));
 sky130_fd_sc_hd__inv_2 _07846_ (.A(_04161_),
    .Y(_04166_));
 sky130_fd_sc_hd__o211a_1 _07847_ (.A1(_04041_),
    .A2(_04166_),
    .B1(_04160_),
    .C1(_04162_),
    .X(_03439_));
 sky130_fd_sc_hd__buf_1 _07848_ (.A(_03991_),
    .X(_04167_));
 sky130_fd_sc_hd__or2_1 _07849_ (.A(_04108_),
    .B(_04033_),
    .X(_04168_));
 sky130_fd_sc_hd__o21ai_1 _07850_ (.A1(_04167_),
    .A2(_04011_),
    .B1(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__inv_2 _07851_ (.A(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__inv_2 _07852_ (.A(_04035_),
    .Y(_04171_));
 sky130_fd_sc_hd__o221a_1 _07853_ (.A1(_04035_),
    .A2(_04170_),
    .B1(_04171_),
    .B2(_04169_),
    .C1(_04165_),
    .X(_03438_));
 sky130_fd_sc_hd__inv_2 _07854_ (.A(_04033_),
    .Y(_04172_));
 sky130_fd_sc_hd__o211a_1 _07855_ (.A1(_04109_),
    .A2(_04172_),
    .B1(_04160_),
    .C1(_04168_),
    .X(_03437_));
 sky130_fd_sc_hd__clkbuf_1 _07856_ (.A(_04106_),
    .X(_04173_));
 sky130_fd_sc_hd__o221a_1 _07857_ (.A1(_03989_),
    .A2(_04042_),
    .B1(_04173_),
    .B2(_04051_),
    .C1(_04043_),
    .X(_04174_));
 sky130_fd_sc_hd__or2_1 _07858_ (.A(_04046_),
    .B(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__o21ai_1 _07859_ (.A1(_04167_),
    .A2(_04044_),
    .B1(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__inv_2 _07860_ (.A(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__inv_2 _07861_ (.A(_04047_),
    .Y(_04178_));
 sky130_fd_sc_hd__o221a_1 _07862_ (.A1(_04047_),
    .A2(_04177_),
    .B1(_04178_),
    .B2(_04176_),
    .C1(_04165_),
    .X(_03436_));
 sky130_fd_sc_hd__nand2_1 _07863_ (.A(_04046_),
    .B(_04174_),
    .Y(_04179_));
 sky130_fd_sc_hd__and3_1 _07864_ (.A(_04153_),
    .B(_04175_),
    .C(_04179_),
    .X(_03435_));
 sky130_fd_sc_hd__or2_1 _07865_ (.A(_04173_),
    .B(_04049_),
    .X(_04180_));
 sky130_fd_sc_hd__o21ai_2 _07866_ (.A1(_04167_),
    .A2(_04042_),
    .B1(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__inv_2 _07867_ (.A(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__inv_2 _07868_ (.A(_04050_),
    .Y(_04183_));
 sky130_fd_sc_hd__buf_1 _07869_ (.A(_04138_),
    .X(_04184_));
 sky130_fd_sc_hd__o221a_1 _07870_ (.A1(_04050_),
    .A2(_04182_),
    .B1(_04183_),
    .B2(_04181_),
    .C1(_04184_),
    .X(_03434_));
 sky130_fd_sc_hd__nand2_1 _07871_ (.A(_04173_),
    .B(_04049_),
    .Y(_04185_));
 sky130_fd_sc_hd__and3_1 _07872_ (.A(_04153_),
    .B(_04180_),
    .C(_04185_),
    .X(_03433_));
 sky130_fd_sc_hd__inv_2 _07873_ (.A(_04059_),
    .Y(_04186_));
 sky130_fd_sc_hd__buf_1 _07874_ (.A(_04068_),
    .X(_04187_));
 sky130_fd_sc_hd__buf_1 _07875_ (.A(_04069_),
    .X(_04188_));
 sky130_fd_sc_hd__buf_1 _07876_ (.A(_04104_),
    .X(_04189_));
 sky130_fd_sc_hd__a31o_1 _07877_ (.A1(_04187_),
    .A2(_04188_),
    .A3(_04189_),
    .B1(_04065_),
    .X(_04190_));
 sky130_fd_sc_hd__nand2_1 _07878_ (.A(_04186_),
    .B(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__o21ai_1 _07879_ (.A1(_04056_),
    .A2(_04058_),
    .B1(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__inv_2 _07880_ (.A(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__o221a_1 _07881_ (.A1(_04055_),
    .A2(_04193_),
    .B1(_04054_),
    .B2(_04192_),
    .C1(_04184_),
    .X(_03432_));
 sky130_fd_sc_hd__buf_1 _07882_ (.A(_03668_),
    .X(_04194_));
 sky130_fd_sc_hd__o211a_1 _07883_ (.A1(_04186_),
    .A2(_04190_),
    .B1(_04194_),
    .C1(_04191_),
    .X(_03431_));
 sky130_fd_sc_hd__nand2_1 _07884_ (.A(_04189_),
    .B(_04188_),
    .Y(_04195_));
 sky130_fd_sc_hd__inv_2 _07885_ (.A(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__o21ai_1 _07886_ (.A1(_04064_),
    .A2(_04196_),
    .B1(_04187_),
    .Y(_04197_));
 sky130_fd_sc_hd__o311a_1 _07887_ (.A1(_04064_),
    .A2(_04196_),
    .A3(_04187_),
    .B1(_03674_),
    .C1(_04197_),
    .X(_03430_));
 sky130_fd_sc_hd__o211a_1 _07888_ (.A1(_04189_),
    .A2(_04188_),
    .B1(_04194_),
    .C1(_04195_),
    .X(_03429_));
 sky130_fd_sc_hd__nand2_1 _07889_ (.A(_04101_),
    .B(_04077_),
    .Y(_04198_));
 sky130_fd_sc_hd__o21ai_1 _07890_ (.A1(_01223_),
    .A2(_04075_),
    .B1(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_1 _07891_ (.A(_04074_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__o211a_1 _07892_ (.A1(_04074_),
    .A2(_04199_),
    .B1(_04194_),
    .C1(_04200_),
    .X(_03428_));
 sky130_fd_sc_hd__buf_1 _07893_ (.A(_03668_),
    .X(_04201_));
 sky130_fd_sc_hd__o211a_1 _07894_ (.A1(_04101_),
    .A2(_04077_),
    .B1(_04201_),
    .C1(_04198_),
    .X(_03427_));
 sky130_fd_sc_hd__or2_1 _07895_ (.A(_04097_),
    .B(_04084_),
    .X(_04202_));
 sky130_fd_sc_hd__o21ai_1 _07896_ (.A1(_04081_),
    .A2(_04083_),
    .B1(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__nand2_1 _07897_ (.A(_04080_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__o211a_1 _07898_ (.A1(_04080_),
    .A2(_04203_),
    .B1(_04201_),
    .C1(_04204_),
    .X(_03426_));
 sky130_fd_sc_hd__o211a_1 _07899_ (.A1(_04098_),
    .A2(_04085_),
    .B1(_04201_),
    .C1(_04202_),
    .X(_03425_));
 sky130_fd_sc_hd__inv_2 _07900_ (.A(_04096_),
    .Y(_04205_));
 sky130_fd_sc_hd__a21oi_2 _07901_ (.A1(_04086_),
    .A2(\e1.offset[3] ),
    .B1(_04087_),
    .Y(_04206_));
 sky130_fd_sc_hd__inv_2 _07902_ (.A(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__o221a_1 _07903_ (.A1(_04205_),
    .A2(_04206_),
    .B1(_04096_),
    .B2(_04207_),
    .C1(_04184_),
    .X(_03424_));
 sky130_fd_sc_hd__a21oi_2 _07904_ (.A1(_04088_),
    .A2(\e1.offset[2] ),
    .B1(_04089_),
    .Y(_04208_));
 sky130_fd_sc_hd__inv_2 _07905_ (.A(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__o221a_1 _07906_ (.A1(_04094_),
    .A2(_04208_),
    .B1(_04095_),
    .B2(_04209_),
    .C1(_04158_),
    .X(_03423_));
 sky130_fd_sc_hd__buf_1 _07907_ (.A(_01211_),
    .X(_04210_));
 sky130_fd_sc_hd__o21a_1 _07908_ (.A1(_04210_),
    .A2(_04091_),
    .B1(_04092_),
    .X(_04211_));
 sky130_fd_sc_hd__and3b_1 _07909_ (.A_N(_04211_),
    .B(_04093_),
    .C(_03669_),
    .X(_03422_));
 sky130_fd_sc_hd__inv_2 _07910_ (.A(_04210_),
    .Y(_04212_));
 sky130_fd_sc_hd__o221a_1 _07911_ (.A1(_04210_),
    .A2(_04091_),
    .B1(_04212_),
    .B2(\e1.offset[0] ),
    .C1(_04158_),
    .X(_03421_));
 sky130_fd_sc_hd__clkbuf_1 _07912_ (.A(_02396_),
    .X(_02395_));
 sky130_fd_sc_hd__clkbuf_1 _07913_ (.A(\r1.waddr[4] ),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _07914_ (.A(\r1.waddr[3] ),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_1 _07915_ (.A(\r1.waddr[2] ),
    .X(_04215_));
 sky130_fd_sc_hd__or3_1 _07916_ (.A(_04213_),
    .B(_04214_),
    .C(_04215_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _07917_ (.A(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__inv_2 _07918_ (.A(\r1.waddr[1] ),
    .Y(_04218_));
 sky130_fd_sc_hd__inv_2 _07919_ (.A(\w1.instruction[5] ),
    .Y(_04219_));
 sky130_fd_sc_hd__o211ai_1 _07920_ (.A1(_04219_),
    .A2(\w1.instruction[4] ),
    .B1(\w1.instruction[1] ),
    .C1(\w1.instruction[0] ),
    .Y(_04220_));
 sky130_fd_sc_hd__or4_4 _07921_ (.A(\w1.instruction[3] ),
    .B(\w1.instruction[2] ),
    .C(\w1.instruction[6] ),
    .D(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__or2b_1 _07922_ (.A(_04221_),
    .B_N(\r1.waddr[0] ),
    .X(_04222_));
 sky130_fd_sc_hd__or2_1 _07923_ (.A(_04218_),
    .B(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__buf_1 _07924_ (.A(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__or2_2 _07925_ (.A(_04217_),
    .B(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__buf_1 _07926_ (.A(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__buf_1 _07927_ (.A(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__buf_1 _07928_ (.A(\r1.wdata[31] ),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_2 _07929_ (.A(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__inv_2 _07930_ (.A(_04225_),
    .Y(_04230_));
 sky130_fd_sc_hd__buf_1 _07931_ (.A(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__buf_1 _07932_ (.A(_04231_),
    .X(_04232_));
 sky130_fd_sc_hd__a22o_1 _07933_ (.A1(\r1.regblock[3][31] ),
    .A2(_04227_),
    .B1(_04229_),
    .B2(_04232_),
    .X(_03420_));
 sky130_fd_sc_hd__clkbuf_1 _07934_ (.A(_02396_),
    .X(_02394_));
 sky130_fd_sc_hd__buf_1 _07935_ (.A(\r1.wdata[30] ),
    .X(_04233_));
 sky130_fd_sc_hd__buf_1 _07936_ (.A(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__a22o_1 _07937_ (.A1(\r1.regblock[3][30] ),
    .A2(_04227_),
    .B1(_04234_),
    .B2(_04232_),
    .X(_03419_));
 sky130_fd_sc_hd__clkbuf_1 _07938_ (.A(_03908_),
    .X(_04235_));
 sky130_fd_sc_hd__buf_2 _07939_ (.A(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_2 _07940_ (.A(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__buf_1 _07941_ (.A(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__buf_1 _07942_ (.A(_04238_),
    .X(_02393_));
 sky130_fd_sc_hd__buf_1 _07943_ (.A(\r1.wdata[29] ),
    .X(_04239_));
 sky130_fd_sc_hd__buf_1 _07944_ (.A(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__a22o_1 _07945_ (.A1(\r1.regblock[3][29] ),
    .A2(_04227_),
    .B1(_04240_),
    .B2(_04232_),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _07946_ (.A(_04238_),
    .X(_02392_));
 sky130_fd_sc_hd__clkbuf_4 _07947_ (.A(_04225_),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_2 _07948_ (.A(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__buf_1 _07949_ (.A(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__buf_1 _07950_ (.A(\r1.wdata[28] ),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_2 _07951_ (.A(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_4 _07952_ (.A(_04230_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_2 _07953_ (.A(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__buf_1 _07954_ (.A(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__a22o_1 _07955_ (.A1(\r1.regblock[3][28] ),
    .A2(_04243_),
    .B1(_04245_),
    .B2(_04248_),
    .X(_03417_));
 sky130_fd_sc_hd__clkbuf_1 _07956_ (.A(_04238_),
    .X(_02391_));
 sky130_fd_sc_hd__buf_1 _07957_ (.A(\r1.wdata[27] ),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_2 _07958_ (.A(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__a22o_1 _07959_ (.A1(\r1.regblock[3][27] ),
    .A2(_04243_),
    .B1(_04250_),
    .B2(_04248_),
    .X(_03416_));
 sky130_fd_sc_hd__buf_1 _07960_ (.A(_04237_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _07961_ (.A(_04251_),
    .X(_02390_));
 sky130_fd_sc_hd__buf_1 _07962_ (.A(\r1.wdata[26] ),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_2 _07963_ (.A(_04252_),
    .X(_04253_));
 sky130_fd_sc_hd__a22o_1 _07964_ (.A1(\r1.regblock[3][26] ),
    .A2(_04243_),
    .B1(_04253_),
    .B2(_04248_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_1 _07965_ (.A(_04251_),
    .X(_02389_));
 sky130_fd_sc_hd__buf_1 _07966_ (.A(_04242_),
    .X(_04254_));
 sky130_fd_sc_hd__buf_1 _07967_ (.A(\r1.wdata[25] ),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_2 _07968_ (.A(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__buf_1 _07969_ (.A(_04247_),
    .X(_04257_));
 sky130_fd_sc_hd__a22o_1 _07970_ (.A1(\r1.regblock[3][25] ),
    .A2(_04254_),
    .B1(_04256_),
    .B2(_04257_),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _07971_ (.A(_04251_),
    .X(_02388_));
 sky130_fd_sc_hd__buf_1 _07972_ (.A(\r1.wdata[24] ),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_2 _07973_ (.A(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__a22o_1 _07974_ (.A1(\r1.regblock[3][24] ),
    .A2(_04254_),
    .B1(_04259_),
    .B2(_04257_),
    .X(_03413_));
 sky130_fd_sc_hd__buf_1 _07975_ (.A(_04237_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _07976_ (.A(_04260_),
    .X(_02387_));
 sky130_fd_sc_hd__buf_1 _07977_ (.A(\r1.wdata[23] ),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_2 _07978_ (.A(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__a22o_1 _07979_ (.A1(\r1.regblock[3][23] ),
    .A2(_04254_),
    .B1(_04262_),
    .B2(_04257_),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_1 _07980_ (.A(_04260_),
    .X(_02386_));
 sky130_fd_sc_hd__buf_1 _07981_ (.A(_04242_),
    .X(_04263_));
 sky130_fd_sc_hd__buf_1 _07982_ (.A(\r1.wdata[22] ),
    .X(_04264_));
 sky130_fd_sc_hd__buf_1 _07983_ (.A(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__buf_1 _07984_ (.A(_04247_),
    .X(_04266_));
 sky130_fd_sc_hd__a22o_1 _07985_ (.A1(\r1.regblock[3][22] ),
    .A2(_04263_),
    .B1(_04265_),
    .B2(_04266_),
    .X(_03411_));
 sky130_fd_sc_hd__clkbuf_1 _07986_ (.A(_04260_),
    .X(_02385_));
 sky130_fd_sc_hd__buf_1 _07987_ (.A(\r1.wdata[21] ),
    .X(_04267_));
 sky130_fd_sc_hd__buf_1 _07988_ (.A(_04267_),
    .X(_04268_));
 sky130_fd_sc_hd__a22o_1 _07989_ (.A1(\r1.regblock[3][21] ),
    .A2(_04263_),
    .B1(_04268_),
    .B2(_04266_),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_2 _07990_ (.A(_04236_),
    .X(_04269_));
 sky130_fd_sc_hd__buf_1 _07991_ (.A(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_2 _07992_ (.A(_04270_),
    .X(_02384_));
 sky130_fd_sc_hd__buf_1 _07993_ (.A(\r1.wdata[20] ),
    .X(_04271_));
 sky130_fd_sc_hd__buf_1 _07994_ (.A(_04271_),
    .X(_04272_));
 sky130_fd_sc_hd__a22o_1 _07995_ (.A1(\r1.regblock[3][20] ),
    .A2(_04263_),
    .B1(_04272_),
    .B2(_04266_),
    .X(_03409_));
 sky130_fd_sc_hd__clkbuf_1 _07996_ (.A(_04270_),
    .X(_02383_));
 sky130_fd_sc_hd__clkbuf_2 _07997_ (.A(_04241_),
    .X(_04273_));
 sky130_fd_sc_hd__buf_1 _07998_ (.A(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__buf_1 _07999_ (.A(\r1.wdata[19] ),
    .X(_04275_));
 sky130_fd_sc_hd__buf_1 _08000_ (.A(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_2 _08001_ (.A(_04246_),
    .X(_04277_));
 sky130_fd_sc_hd__buf_1 _08002_ (.A(_04277_),
    .X(_04278_));
 sky130_fd_sc_hd__a22o_1 _08003_ (.A1(\r1.regblock[3][19] ),
    .A2(_04274_),
    .B1(_04276_),
    .B2(_04278_),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _08004_ (.A(_04270_),
    .X(_02382_));
 sky130_fd_sc_hd__buf_1 _08005_ (.A(\r1.wdata[18] ),
    .X(_04279_));
 sky130_fd_sc_hd__buf_1 _08006_ (.A(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__a22o_1 _08007_ (.A1(\r1.regblock[3][18] ),
    .A2(_04274_),
    .B1(_04280_),
    .B2(_04278_),
    .X(_03407_));
 sky130_fd_sc_hd__buf_1 _08008_ (.A(_04269_),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _08009_ (.A(_04281_),
    .X(_02381_));
 sky130_fd_sc_hd__buf_1 _08010_ (.A(\r1.wdata[17] ),
    .X(_04282_));
 sky130_fd_sc_hd__buf_1 _08011_ (.A(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__a22o_1 _08012_ (.A1(\r1.regblock[3][17] ),
    .A2(_04274_),
    .B1(_04283_),
    .B2(_04278_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_1 _08013_ (.A(_04281_),
    .X(_02380_));
 sky130_fd_sc_hd__buf_1 _08014_ (.A(_04273_),
    .X(_04284_));
 sky130_fd_sc_hd__buf_1 _08015_ (.A(\r1.wdata[16] ),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_2 _08016_ (.A(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__buf_1 _08017_ (.A(_04277_),
    .X(_04287_));
 sky130_fd_sc_hd__a22o_1 _08018_ (.A1(\r1.regblock[3][16] ),
    .A2(_04284_),
    .B1(_04286_),
    .B2(_04287_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_1 _08019_ (.A(_04281_),
    .X(_02379_));
 sky130_fd_sc_hd__buf_1 _08020_ (.A(\r1.wdata[15] ),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_2 _08021_ (.A(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__a22o_1 _08022_ (.A1(\r1.regblock[3][15] ),
    .A2(_04284_),
    .B1(_04289_),
    .B2(_04287_),
    .X(_03404_));
 sky130_fd_sc_hd__buf_1 _08023_ (.A(_04269_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _08024_ (.A(_04290_),
    .X(_02378_));
 sky130_fd_sc_hd__buf_1 _08025_ (.A(\r1.wdata[14] ),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_2 _08026_ (.A(_04291_),
    .X(_04292_));
 sky130_fd_sc_hd__a22o_1 _08027_ (.A1(\r1.regblock[3][14] ),
    .A2(_04284_),
    .B1(_04292_),
    .B2(_04287_),
    .X(_03403_));
 sky130_fd_sc_hd__clkbuf_1 _08028_ (.A(_04290_),
    .X(_02377_));
 sky130_fd_sc_hd__buf_1 _08029_ (.A(_04273_),
    .X(_04293_));
 sky130_fd_sc_hd__buf_1 _08030_ (.A(\r1.wdata[13] ),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_2 _08031_ (.A(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__buf_1 _08032_ (.A(_04277_),
    .X(_04296_));
 sky130_fd_sc_hd__a22o_1 _08033_ (.A1(\r1.regblock[3][13] ),
    .A2(_04293_),
    .B1(_04295_),
    .B2(_04296_),
    .X(_03402_));
 sky130_fd_sc_hd__clkbuf_1 _08034_ (.A(_04290_),
    .X(_02376_));
 sky130_fd_sc_hd__buf_1 _08035_ (.A(\r1.wdata[12] ),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_2 _08036_ (.A(_04297_),
    .X(_04298_));
 sky130_fd_sc_hd__a22o_1 _08037_ (.A1(\r1.regblock[3][12] ),
    .A2(_04293_),
    .B1(_04298_),
    .B2(_04296_),
    .X(_03401_));
 sky130_fd_sc_hd__buf_1 _08038_ (.A(_04236_),
    .X(_04299_));
 sky130_fd_sc_hd__buf_2 _08039_ (.A(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _08040_ (.A(_04300_),
    .X(_02375_));
 sky130_fd_sc_hd__buf_1 _08041_ (.A(\r1.wdata[11] ),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_2 _08042_ (.A(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__a22o_1 _08043_ (.A1(\r1.regblock[3][11] ),
    .A2(_04293_),
    .B1(_04302_),
    .B2(_04296_),
    .X(_03400_));
 sky130_fd_sc_hd__clkbuf_1 _08044_ (.A(_04300_),
    .X(_02374_));
 sky130_fd_sc_hd__buf_1 _08045_ (.A(_04241_),
    .X(_04303_));
 sky130_fd_sc_hd__buf_1 _08046_ (.A(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__buf_1 _08047_ (.A(\r1.wdata[10] ),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_2 _08048_ (.A(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__buf_1 _08049_ (.A(_04246_),
    .X(_04307_));
 sky130_fd_sc_hd__buf_1 _08050_ (.A(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__a22o_1 _08051_ (.A1(\r1.regblock[3][10] ),
    .A2(_04304_),
    .B1(_04306_),
    .B2(_04308_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_1 _08052_ (.A(_04300_),
    .X(_02373_));
 sky130_fd_sc_hd__buf_1 _08053_ (.A(\r1.wdata[9] ),
    .X(_04309_));
 sky130_fd_sc_hd__clkbuf_2 _08054_ (.A(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__a22o_1 _08055_ (.A1(\r1.regblock[3][9] ),
    .A2(_04304_),
    .B1(_04310_),
    .B2(_04308_),
    .X(_03398_));
 sky130_fd_sc_hd__buf_1 _08056_ (.A(_04299_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _08057_ (.A(_04311_),
    .X(_02372_));
 sky130_fd_sc_hd__buf_1 _08058_ (.A(\r1.wdata[8] ),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_2 _08059_ (.A(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__a22o_1 _08060_ (.A1(\r1.regblock[3][8] ),
    .A2(_04304_),
    .B1(_04313_),
    .B2(_04308_),
    .X(_03397_));
 sky130_fd_sc_hd__clkbuf_1 _08061_ (.A(_04311_),
    .X(_02371_));
 sky130_fd_sc_hd__buf_1 _08062_ (.A(_04303_),
    .X(_04314_));
 sky130_fd_sc_hd__buf_1 _08063_ (.A(\r1.wdata[7] ),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_2 _08064_ (.A(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__buf_1 _08065_ (.A(_04307_),
    .X(_04317_));
 sky130_fd_sc_hd__a22o_1 _08066_ (.A1(\r1.regblock[3][7] ),
    .A2(_04314_),
    .B1(_04316_),
    .B2(_04317_),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_1 _08067_ (.A(_04311_),
    .X(_02370_));
 sky130_fd_sc_hd__buf_1 _08068_ (.A(\r1.wdata[6] ),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_2 _08069_ (.A(_04318_),
    .X(_04319_));
 sky130_fd_sc_hd__a22o_1 _08070_ (.A1(\r1.regblock[3][6] ),
    .A2(_04314_),
    .B1(_04319_),
    .B2(_04317_),
    .X(_03395_));
 sky130_fd_sc_hd__buf_1 _08071_ (.A(_04299_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_1 _08072_ (.A(_04320_),
    .X(_02369_));
 sky130_fd_sc_hd__buf_1 _08073_ (.A(\r1.wdata[5] ),
    .X(_04321_));
 sky130_fd_sc_hd__clkbuf_2 _08074_ (.A(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__a22o_1 _08075_ (.A1(\r1.regblock[3][5] ),
    .A2(_04314_),
    .B1(_04322_),
    .B2(_04317_),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_1 _08076_ (.A(_04320_),
    .X(_02368_));
 sky130_fd_sc_hd__buf_1 _08077_ (.A(_04303_),
    .X(_04323_));
 sky130_fd_sc_hd__buf_1 _08078_ (.A(\r1.wdata[4] ),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_2 _08079_ (.A(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__buf_1 _08080_ (.A(_04307_),
    .X(_04326_));
 sky130_fd_sc_hd__a22o_1 _08081_ (.A1(\r1.regblock[3][4] ),
    .A2(_04323_),
    .B1(_04325_),
    .B2(_04326_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_1 _08082_ (.A(_04320_),
    .X(_02367_));
 sky130_fd_sc_hd__buf_1 _08083_ (.A(\r1.wdata[3] ),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_2 _08084_ (.A(_04327_),
    .X(_04328_));
 sky130_fd_sc_hd__a22o_1 _08085_ (.A1(\r1.regblock[3][3] ),
    .A2(_04323_),
    .B1(_04328_),
    .B2(_04326_),
    .X(_03392_));
 sky130_fd_sc_hd__buf_1 _08086_ (.A(_04235_),
    .X(_04329_));
 sky130_fd_sc_hd__buf_2 _08087_ (.A(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__buf_1 _08088_ (.A(_04330_),
    .X(_04331_));
 sky130_fd_sc_hd__buf_1 _08089_ (.A(_04331_),
    .X(_02366_));
 sky130_fd_sc_hd__buf_1 _08090_ (.A(\r1.wdata[2] ),
    .X(_04332_));
 sky130_fd_sc_hd__clkbuf_2 _08091_ (.A(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__a22o_1 _08092_ (.A1(\r1.regblock[3][2] ),
    .A2(_04323_),
    .B1(_04333_),
    .B2(_04326_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_1 _08093_ (.A(_04331_),
    .X(_02365_));
 sky130_fd_sc_hd__buf_1 _08094_ (.A(\r1.wdata[1] ),
    .X(_04334_));
 sky130_fd_sc_hd__buf_1 _08095_ (.A(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__a22o_1 _08096_ (.A1(\r1.regblock[3][1] ),
    .A2(_04226_),
    .B1(_04335_),
    .B2(_04231_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _08097_ (.A(_04331_),
    .X(_02364_));
 sky130_fd_sc_hd__buf_1 _08098_ (.A(\r1.wdata[0] ),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_2 _08099_ (.A(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__a22o_1 _08100_ (.A1(\r1.regblock[3][0] ),
    .A2(_04226_),
    .B1(_04337_),
    .B2(_04231_),
    .X(_03389_));
 sky130_fd_sc_hd__buf_1 _08101_ (.A(_04330_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _08102_ (.A(_04338_),
    .X(_02363_));
 sky130_fd_sc_hd__clkbuf_1 _08103_ (.A(_04224_),
    .X(_04339_));
 sky130_fd_sc_hd__inv_2 _08104_ (.A(\r1.waddr[4] ),
    .Y(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _08105_ (.A(_04340_),
    .X(_04341_));
 sky130_fd_sc_hd__or3_1 _08106_ (.A(_04341_),
    .B(_04214_),
    .C(_04215_),
    .X(_04342_));
 sky130_fd_sc_hd__or2_2 _08107_ (.A(_04339_),
    .B(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_2 _08108_ (.A(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__buf_1 _08109_ (.A(_04344_),
    .X(_04345_));
 sky130_fd_sc_hd__inv_2 _08110_ (.A(_04343_),
    .Y(_04346_));
 sky130_fd_sc_hd__clkbuf_2 _08111_ (.A(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__buf_1 _08112_ (.A(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__a22o_1 _08113_ (.A1(\r1.regblock[19][31] ),
    .A2(_04345_),
    .B1(_04229_),
    .B2(_04348_),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_1 _08114_ (.A(_04338_),
    .X(_02362_));
 sky130_fd_sc_hd__a22o_1 _08115_ (.A1(\r1.regblock[19][30] ),
    .A2(_04345_),
    .B1(_04234_),
    .B2(_04348_),
    .X(_03387_));
 sky130_fd_sc_hd__clkbuf_1 _08116_ (.A(_04338_),
    .X(_02361_));
 sky130_fd_sc_hd__a22o_1 _08117_ (.A1(\r1.regblock[19][29] ),
    .A2(_04345_),
    .B1(_04240_),
    .B2(_04348_),
    .X(_03386_));
 sky130_fd_sc_hd__buf_1 _08118_ (.A(_04330_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _08119_ (.A(_04349_),
    .X(_02360_));
 sky130_fd_sc_hd__clkbuf_2 _08120_ (.A(_04343_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_4 _08121_ (.A(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__buf_1 _08122_ (.A(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_2 _08123_ (.A(_04346_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_4 _08124_ (.A(_04353_),
    .X(_04354_));
 sky130_fd_sc_hd__buf_1 _08125_ (.A(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__a22o_1 _08126_ (.A1(\r1.regblock[19][28] ),
    .A2(_04352_),
    .B1(_04245_),
    .B2(_04355_),
    .X(_03385_));
 sky130_fd_sc_hd__clkbuf_1 _08127_ (.A(_04349_),
    .X(_02359_));
 sky130_fd_sc_hd__a22o_1 _08128_ (.A1(\r1.regblock[19][27] ),
    .A2(_04352_),
    .B1(_04250_),
    .B2(_04355_),
    .X(_03384_));
 sky130_fd_sc_hd__clkbuf_1 _08129_ (.A(_04349_),
    .X(_02358_));
 sky130_fd_sc_hd__a22o_1 _08130_ (.A1(\r1.regblock[19][26] ),
    .A2(_04352_),
    .B1(_04253_),
    .B2(_04355_),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_4 _08131_ (.A(_04329_),
    .X(_04356_));
 sky130_fd_sc_hd__buf_1 _08132_ (.A(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _08133_ (.A(_04357_),
    .X(_02357_));
 sky130_fd_sc_hd__buf_1 _08134_ (.A(_04351_),
    .X(_04358_));
 sky130_fd_sc_hd__buf_1 _08135_ (.A(_04354_),
    .X(_04359_));
 sky130_fd_sc_hd__a22o_1 _08136_ (.A1(\r1.regblock[19][25] ),
    .A2(_04358_),
    .B1(_04256_),
    .B2(_04359_),
    .X(_03382_));
 sky130_fd_sc_hd__clkbuf_1 _08137_ (.A(_04357_),
    .X(_02356_));
 sky130_fd_sc_hd__a22o_1 _08138_ (.A1(\r1.regblock[19][24] ),
    .A2(_04358_),
    .B1(_04259_),
    .B2(_04359_),
    .X(_03381_));
 sky130_fd_sc_hd__clkbuf_1 _08139_ (.A(_04357_),
    .X(_02355_));
 sky130_fd_sc_hd__a22o_1 _08140_ (.A1(\r1.regblock[19][23] ),
    .A2(_04358_),
    .B1(_04262_),
    .B2(_04359_),
    .X(_03380_));
 sky130_fd_sc_hd__buf_1 _08141_ (.A(_04356_),
    .X(_04360_));
 sky130_fd_sc_hd__clkbuf_1 _08142_ (.A(_04360_),
    .X(_02354_));
 sky130_fd_sc_hd__buf_1 _08143_ (.A(_04351_),
    .X(_04361_));
 sky130_fd_sc_hd__buf_1 _08144_ (.A(_04354_),
    .X(_04362_));
 sky130_fd_sc_hd__a22o_1 _08145_ (.A1(\r1.regblock[19][22] ),
    .A2(_04361_),
    .B1(_04265_),
    .B2(_04362_),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_1 _08146_ (.A(_04360_),
    .X(_02353_));
 sky130_fd_sc_hd__a22o_1 _08147_ (.A1(\r1.regblock[19][21] ),
    .A2(_04361_),
    .B1(_04268_),
    .B2(_04362_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_1 _08148_ (.A(_04360_),
    .X(_02352_));
 sky130_fd_sc_hd__a22o_1 _08149_ (.A1(\r1.regblock[19][20] ),
    .A2(_04361_),
    .B1(_04272_),
    .B2(_04362_),
    .X(_03377_));
 sky130_fd_sc_hd__buf_1 _08150_ (.A(_04356_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _08151_ (.A(_04363_),
    .X(_02351_));
 sky130_fd_sc_hd__buf_2 _08152_ (.A(_04350_),
    .X(_04364_));
 sky130_fd_sc_hd__buf_1 _08153_ (.A(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__buf_2 _08154_ (.A(_04353_),
    .X(_04366_));
 sky130_fd_sc_hd__buf_1 _08155_ (.A(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__a22o_1 _08156_ (.A1(\r1.regblock[19][19] ),
    .A2(_04365_),
    .B1(_04276_),
    .B2(_04367_),
    .X(_03376_));
 sky130_fd_sc_hd__clkbuf_1 _08157_ (.A(_04363_),
    .X(_02350_));
 sky130_fd_sc_hd__a22o_1 _08158_ (.A1(\r1.regblock[19][18] ),
    .A2(_04365_),
    .B1(_04280_),
    .B2(_04367_),
    .X(_03375_));
 sky130_fd_sc_hd__clkbuf_1 _08159_ (.A(_04363_),
    .X(_02349_));
 sky130_fd_sc_hd__a22o_1 _08160_ (.A1(\r1.regblock[19][17] ),
    .A2(_04365_),
    .B1(_04283_),
    .B2(_04367_),
    .X(_03374_));
 sky130_fd_sc_hd__buf_4 _08161_ (.A(_04329_),
    .X(_04368_));
 sky130_fd_sc_hd__clkbuf_1 _08162_ (.A(_04368_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _08163_ (.A(_04369_),
    .X(_02348_));
 sky130_fd_sc_hd__buf_1 _08164_ (.A(_04364_),
    .X(_04370_));
 sky130_fd_sc_hd__buf_1 _08165_ (.A(_04366_),
    .X(_04371_));
 sky130_fd_sc_hd__a22o_1 _08166_ (.A1(\r1.regblock[19][16] ),
    .A2(_04370_),
    .B1(_04286_),
    .B2(_04371_),
    .X(_03373_));
 sky130_fd_sc_hd__clkbuf_1 _08167_ (.A(_04369_),
    .X(_02347_));
 sky130_fd_sc_hd__a22o_1 _08168_ (.A1(\r1.regblock[19][15] ),
    .A2(_04370_),
    .B1(_04289_),
    .B2(_04371_),
    .X(_03372_));
 sky130_fd_sc_hd__clkbuf_1 _08169_ (.A(_04369_),
    .X(_02346_));
 sky130_fd_sc_hd__a22o_1 _08170_ (.A1(\r1.regblock[19][14] ),
    .A2(_04370_),
    .B1(_04292_),
    .B2(_04371_),
    .X(_03371_));
 sky130_fd_sc_hd__buf_1 _08171_ (.A(_04368_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _08172_ (.A(_04372_),
    .X(_02345_));
 sky130_fd_sc_hd__buf_1 _08173_ (.A(_04364_),
    .X(_04373_));
 sky130_fd_sc_hd__buf_1 _08174_ (.A(_04366_),
    .X(_04374_));
 sky130_fd_sc_hd__a22o_1 _08175_ (.A1(\r1.regblock[19][13] ),
    .A2(_04373_),
    .B1(_04295_),
    .B2(_04374_),
    .X(_03370_));
 sky130_fd_sc_hd__clkbuf_1 _08176_ (.A(_04372_),
    .X(_02344_));
 sky130_fd_sc_hd__a22o_1 _08177_ (.A1(\r1.regblock[19][12] ),
    .A2(_04373_),
    .B1(_04298_),
    .B2(_04374_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_1 _08178_ (.A(_04372_),
    .X(_02343_));
 sky130_fd_sc_hd__a22o_1 _08179_ (.A1(\r1.regblock[19][11] ),
    .A2(_04373_),
    .B1(_04302_),
    .B2(_04374_),
    .X(_03368_));
 sky130_fd_sc_hd__buf_1 _08180_ (.A(_04368_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_1 _08181_ (.A(_04375_),
    .X(_02342_));
 sky130_fd_sc_hd__clkbuf_2 _08182_ (.A(_04350_),
    .X(_04376_));
 sky130_fd_sc_hd__buf_1 _08183_ (.A(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_2 _08184_ (.A(_04353_),
    .X(_04378_));
 sky130_fd_sc_hd__buf_1 _08185_ (.A(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__a22o_1 _08186_ (.A1(\r1.regblock[19][10] ),
    .A2(_04377_),
    .B1(_04306_),
    .B2(_04379_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_1 _08187_ (.A(_04375_),
    .X(_02341_));
 sky130_fd_sc_hd__a22o_1 _08188_ (.A1(\r1.regblock[19][9] ),
    .A2(_04377_),
    .B1(_04310_),
    .B2(_04379_),
    .X(_03366_));
 sky130_fd_sc_hd__clkbuf_1 _08189_ (.A(_04375_),
    .X(_02340_));
 sky130_fd_sc_hd__a22o_1 _08190_ (.A1(\r1.regblock[19][8] ),
    .A2(_04377_),
    .B1(_04313_),
    .B2(_04379_),
    .X(_03365_));
 sky130_fd_sc_hd__clkbuf_2 _08191_ (.A(_04235_),
    .X(_04380_));
 sky130_fd_sc_hd__buf_1 _08192_ (.A(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__buf_1 _08193_ (.A(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _08194_ (.A(_04382_),
    .X(_02339_));
 sky130_fd_sc_hd__buf_1 _08195_ (.A(_04376_),
    .X(_04383_));
 sky130_fd_sc_hd__buf_1 _08196_ (.A(_04378_),
    .X(_04384_));
 sky130_fd_sc_hd__a22o_1 _08197_ (.A1(\r1.regblock[19][7] ),
    .A2(_04383_),
    .B1(_04316_),
    .B2(_04384_),
    .X(_03364_));
 sky130_fd_sc_hd__clkbuf_1 _08198_ (.A(_04382_),
    .X(_02338_));
 sky130_fd_sc_hd__a22o_1 _08199_ (.A1(\r1.regblock[19][6] ),
    .A2(_04383_),
    .B1(_04319_),
    .B2(_04384_),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_1 _08200_ (.A(_04382_),
    .X(_02337_));
 sky130_fd_sc_hd__a22o_1 _08201_ (.A1(\r1.regblock[19][5] ),
    .A2(_04383_),
    .B1(_04322_),
    .B2(_04384_),
    .X(_03362_));
 sky130_fd_sc_hd__buf_1 _08202_ (.A(_04381_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _08203_ (.A(_04385_),
    .X(_02336_));
 sky130_fd_sc_hd__buf_1 _08204_ (.A(_04376_),
    .X(_04386_));
 sky130_fd_sc_hd__buf_1 _08205_ (.A(_04378_),
    .X(_04387_));
 sky130_fd_sc_hd__a22o_1 _08206_ (.A1(\r1.regblock[19][4] ),
    .A2(_04386_),
    .B1(_04325_),
    .B2(_04387_),
    .X(_03361_));
 sky130_fd_sc_hd__clkbuf_1 _08207_ (.A(_04385_),
    .X(_02335_));
 sky130_fd_sc_hd__a22o_1 _08208_ (.A1(\r1.regblock[19][3] ),
    .A2(_04386_),
    .B1(_04328_),
    .B2(_04387_),
    .X(_03360_));
 sky130_fd_sc_hd__clkbuf_1 _08209_ (.A(_04385_),
    .X(_02334_));
 sky130_fd_sc_hd__a22o_1 _08210_ (.A1(\r1.regblock[19][2] ),
    .A2(_04386_),
    .B1(_04333_),
    .B2(_04387_),
    .X(_03359_));
 sky130_fd_sc_hd__clkbuf_2 _08211_ (.A(_04381_),
    .X(_04388_));
 sky130_fd_sc_hd__clkbuf_1 _08212_ (.A(_04388_),
    .X(_02333_));
 sky130_fd_sc_hd__a22o_1 _08213_ (.A1(\r1.regblock[19][1] ),
    .A2(_04344_),
    .B1(_04335_),
    .B2(_04347_),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_1 _08214_ (.A(_04388_),
    .X(_02332_));
 sky130_fd_sc_hd__a22o_1 _08215_ (.A1(\r1.regblock[19][0] ),
    .A2(_04344_),
    .B1(_04337_),
    .B2(_04347_),
    .X(_03357_));
 sky130_fd_sc_hd__clkbuf_1 _08216_ (.A(_04388_),
    .X(_02331_));
 sky130_fd_sc_hd__inv_2 _08217_ (.A(\r1.waddr[3] ),
    .Y(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _08218_ (.A(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__inv_2 _08219_ (.A(\r1.waddr[2] ),
    .Y(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _08220_ (.A(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__or3_1 _08221_ (.A(_04213_),
    .B(_04390_),
    .C(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__clkbuf_1 _08222_ (.A(_04393_),
    .X(_04394_));
 sky130_fd_sc_hd__or2_1 _08223_ (.A(\r1.waddr[1] ),
    .B(_04222_),
    .X(_04395_));
 sky130_fd_sc_hd__buf_1 _08224_ (.A(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__or2_2 _08225_ (.A(_04394_),
    .B(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__buf_1 _08226_ (.A(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__buf_1 _08227_ (.A(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__inv_2 _08228_ (.A(_04397_),
    .Y(_04400_));
 sky130_fd_sc_hd__buf_1 _08229_ (.A(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__buf_1 _08230_ (.A(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__a22o_1 _08231_ (.A1(\r1.regblock[13][31] ),
    .A2(_04399_),
    .B1(_04229_),
    .B2(_04402_),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_4 _08232_ (.A(_04380_),
    .X(_04403_));
 sky130_fd_sc_hd__buf_1 _08233_ (.A(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__clkbuf_1 _08234_ (.A(_04404_),
    .X(_02330_));
 sky130_fd_sc_hd__a22o_1 _08235_ (.A1(\r1.regblock[13][30] ),
    .A2(_04399_),
    .B1(_04234_),
    .B2(_04402_),
    .X(_03355_));
 sky130_fd_sc_hd__clkbuf_1 _08236_ (.A(_04404_),
    .X(_02329_));
 sky130_fd_sc_hd__a22o_1 _08237_ (.A1(\r1.regblock[13][29] ),
    .A2(_04399_),
    .B1(_04240_),
    .B2(_04402_),
    .X(_03354_));
 sky130_fd_sc_hd__buf_1 _08238_ (.A(_04404_),
    .X(_02328_));
 sky130_fd_sc_hd__clkbuf_4 _08239_ (.A(_04397_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_2 _08240_ (.A(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__buf_1 _08241_ (.A(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_4 _08242_ (.A(_04400_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_2 _08243_ (.A(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__buf_1 _08244_ (.A(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__a22o_1 _08245_ (.A1(\r1.regblock[13][28] ),
    .A2(_04407_),
    .B1(_04245_),
    .B2(_04410_),
    .X(_03353_));
 sky130_fd_sc_hd__buf_1 _08246_ (.A(_04403_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _08247_ (.A(_04411_),
    .X(_02327_));
 sky130_fd_sc_hd__a22o_1 _08248_ (.A1(\r1.regblock[13][27] ),
    .A2(_04407_),
    .B1(_04250_),
    .B2(_04410_),
    .X(_03352_));
 sky130_fd_sc_hd__clkbuf_1 _08249_ (.A(_04411_),
    .X(_02326_));
 sky130_fd_sc_hd__a22o_1 _08250_ (.A1(\r1.regblock[13][26] ),
    .A2(_04407_),
    .B1(_04253_),
    .B2(_04410_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_1 _08251_ (.A(_04411_),
    .X(_02325_));
 sky130_fd_sc_hd__buf_1 _08252_ (.A(_04406_),
    .X(_04412_));
 sky130_fd_sc_hd__buf_1 _08253_ (.A(_04409_),
    .X(_04413_));
 sky130_fd_sc_hd__a22o_1 _08254_ (.A1(\r1.regblock[13][25] ),
    .A2(_04412_),
    .B1(_04256_),
    .B2(_04413_),
    .X(_03350_));
 sky130_fd_sc_hd__buf_1 _08255_ (.A(_04403_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_1 _08256_ (.A(_04414_),
    .X(_02324_));
 sky130_fd_sc_hd__a22o_1 _08257_ (.A1(\r1.regblock[13][24] ),
    .A2(_04412_),
    .B1(_04259_),
    .B2(_04413_),
    .X(_03349_));
 sky130_fd_sc_hd__clkbuf_1 _08258_ (.A(_04414_),
    .X(_02323_));
 sky130_fd_sc_hd__a22o_1 _08259_ (.A1(\r1.regblock[13][23] ),
    .A2(_04412_),
    .B1(_04262_),
    .B2(_04413_),
    .X(_03348_));
 sky130_fd_sc_hd__clkbuf_1 _08260_ (.A(_04414_),
    .X(_02322_));
 sky130_fd_sc_hd__buf_1 _08261_ (.A(_04406_),
    .X(_04415_));
 sky130_fd_sc_hd__buf_1 _08262_ (.A(_04409_),
    .X(_04416_));
 sky130_fd_sc_hd__a22o_1 _08263_ (.A1(\r1.regblock[13][22] ),
    .A2(_04415_),
    .B1(_04265_),
    .B2(_04416_),
    .X(_03347_));
 sky130_fd_sc_hd__buf_1 _08264_ (.A(_04380_),
    .X(_04417_));
 sky130_fd_sc_hd__buf_2 _08265_ (.A(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_1 _08266_ (.A(_04418_),
    .X(_02321_));
 sky130_fd_sc_hd__a22o_1 _08267_ (.A1(\r1.regblock[13][21] ),
    .A2(_04415_),
    .B1(_04268_),
    .B2(_04416_),
    .X(_03346_));
 sky130_fd_sc_hd__clkbuf_1 _08268_ (.A(_04418_),
    .X(_02320_));
 sky130_fd_sc_hd__a22o_1 _08269_ (.A1(\r1.regblock[13][20] ),
    .A2(_04415_),
    .B1(_04272_),
    .B2(_04416_),
    .X(_03345_));
 sky130_fd_sc_hd__clkbuf_1 _08270_ (.A(_04418_),
    .X(_02319_));
 sky130_fd_sc_hd__clkbuf_2 _08271_ (.A(_04405_),
    .X(_04419_));
 sky130_fd_sc_hd__buf_1 _08272_ (.A(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__clkbuf_2 _08273_ (.A(_04408_),
    .X(_04421_));
 sky130_fd_sc_hd__buf_1 _08274_ (.A(_04421_),
    .X(_04422_));
 sky130_fd_sc_hd__a22o_1 _08275_ (.A1(\r1.regblock[13][19] ),
    .A2(_04420_),
    .B1(_04276_),
    .B2(_04422_),
    .X(_03344_));
 sky130_fd_sc_hd__buf_1 _08276_ (.A(_04417_),
    .X(_04423_));
 sky130_fd_sc_hd__clkbuf_1 _08277_ (.A(_04423_),
    .X(_02318_));
 sky130_fd_sc_hd__a22o_1 _08278_ (.A1(\r1.regblock[13][18] ),
    .A2(_04420_),
    .B1(_04280_),
    .B2(_04422_),
    .X(_03343_));
 sky130_fd_sc_hd__clkbuf_1 _08279_ (.A(_04423_),
    .X(_02317_));
 sky130_fd_sc_hd__a22o_1 _08280_ (.A1(\r1.regblock[13][17] ),
    .A2(_04420_),
    .B1(_04283_),
    .B2(_04422_),
    .X(_03342_));
 sky130_fd_sc_hd__clkbuf_1 _08281_ (.A(_04423_),
    .X(_02316_));
 sky130_fd_sc_hd__buf_1 _08282_ (.A(_04419_),
    .X(_04424_));
 sky130_fd_sc_hd__buf_1 _08283_ (.A(_04421_),
    .X(_04425_));
 sky130_fd_sc_hd__a22o_1 _08284_ (.A1(\r1.regblock[13][16] ),
    .A2(_04424_),
    .B1(_04286_),
    .B2(_04425_),
    .X(_03341_));
 sky130_fd_sc_hd__buf_1 _08285_ (.A(_04417_),
    .X(_04426_));
 sky130_fd_sc_hd__clkbuf_1 _08286_ (.A(_04426_),
    .X(_02315_));
 sky130_fd_sc_hd__a22o_1 _08287_ (.A1(\r1.regblock[13][15] ),
    .A2(_04424_),
    .B1(_04289_),
    .B2(_04425_),
    .X(_03340_));
 sky130_fd_sc_hd__clkbuf_1 _08288_ (.A(_04426_),
    .X(_02314_));
 sky130_fd_sc_hd__a22o_1 _08289_ (.A1(\r1.regblock[13][14] ),
    .A2(_04424_),
    .B1(_04292_),
    .B2(_04425_),
    .X(_03339_));
 sky130_fd_sc_hd__clkbuf_1 _08290_ (.A(_04426_),
    .X(_02313_));
 sky130_fd_sc_hd__buf_1 _08291_ (.A(_04419_),
    .X(_04427_));
 sky130_fd_sc_hd__buf_1 _08292_ (.A(_04421_),
    .X(_04428_));
 sky130_fd_sc_hd__a22o_1 _08293_ (.A1(\r1.regblock[13][13] ),
    .A2(_04427_),
    .B1(_04295_),
    .B2(_04428_),
    .X(_03338_));
 sky130_fd_sc_hd__buf_1 _08294_ (.A(net55),
    .X(_04429_));
 sky130_fd_sc_hd__buf_1 _08295_ (.A(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_1 _08296_ (.A(_04430_),
    .X(_04431_));
 sky130_fd_sc_hd__buf_2 _08297_ (.A(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__buf_1 _08298_ (.A(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__buf_2 _08299_ (.A(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__clkbuf_1 _08300_ (.A(_04434_),
    .X(_02312_));
 sky130_fd_sc_hd__a22o_1 _08301_ (.A1(\r1.regblock[13][12] ),
    .A2(_04427_),
    .B1(_04298_),
    .B2(_04428_),
    .X(_03337_));
 sky130_fd_sc_hd__clkbuf_1 _08302_ (.A(_04434_),
    .X(_02311_));
 sky130_fd_sc_hd__a22o_1 _08303_ (.A1(\r1.regblock[13][11] ),
    .A2(_04427_),
    .B1(_04302_),
    .B2(_04428_),
    .X(_03336_));
 sky130_fd_sc_hd__clkbuf_1 _08304_ (.A(_04434_),
    .X(_02310_));
 sky130_fd_sc_hd__buf_1 _08305_ (.A(_04405_),
    .X(_04435_));
 sky130_fd_sc_hd__buf_1 _08306_ (.A(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__buf_1 _08307_ (.A(_04408_),
    .X(_04437_));
 sky130_fd_sc_hd__buf_1 _08308_ (.A(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__a22o_1 _08309_ (.A1(\r1.regblock[13][10] ),
    .A2(_04436_),
    .B1(_04306_),
    .B2(_04438_),
    .X(_03335_));
 sky130_fd_sc_hd__buf_1 _08310_ (.A(_04433_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _08311_ (.A(_04439_),
    .X(_02309_));
 sky130_fd_sc_hd__a22o_1 _08312_ (.A1(\r1.regblock[13][9] ),
    .A2(_04436_),
    .B1(_04310_),
    .B2(_04438_),
    .X(_03334_));
 sky130_fd_sc_hd__clkbuf_1 _08313_ (.A(_04439_),
    .X(_02308_));
 sky130_fd_sc_hd__a22o_1 _08314_ (.A1(\r1.regblock[13][8] ),
    .A2(_04436_),
    .B1(_04313_),
    .B2(_04438_),
    .X(_03333_));
 sky130_fd_sc_hd__clkbuf_1 _08315_ (.A(_04439_),
    .X(_02307_));
 sky130_fd_sc_hd__buf_1 _08316_ (.A(_04435_),
    .X(_04440_));
 sky130_fd_sc_hd__buf_1 _08317_ (.A(_04437_),
    .X(_04441_));
 sky130_fd_sc_hd__a22o_1 _08318_ (.A1(\r1.regblock[13][7] ),
    .A2(_04440_),
    .B1(_04316_),
    .B2(_04441_),
    .X(_03332_));
 sky130_fd_sc_hd__buf_1 _08319_ (.A(_04433_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_1 _08320_ (.A(_04442_),
    .X(_02306_));
 sky130_fd_sc_hd__a22o_1 _08321_ (.A1(\r1.regblock[13][6] ),
    .A2(_04440_),
    .B1(_04319_),
    .B2(_04441_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_1 _08322_ (.A(_04442_),
    .X(_02305_));
 sky130_fd_sc_hd__a22o_1 _08323_ (.A1(\r1.regblock[13][5] ),
    .A2(_04440_),
    .B1(_04322_),
    .B2(_04441_),
    .X(_03330_));
 sky130_fd_sc_hd__clkbuf_1 _08324_ (.A(_04442_),
    .X(_02304_));
 sky130_fd_sc_hd__buf_1 _08325_ (.A(_04435_),
    .X(_04443_));
 sky130_fd_sc_hd__buf_1 _08326_ (.A(_04437_),
    .X(_04444_));
 sky130_fd_sc_hd__a22o_1 _08327_ (.A1(\r1.regblock[13][4] ),
    .A2(_04443_),
    .B1(_04325_),
    .B2(_04444_),
    .X(_03329_));
 sky130_fd_sc_hd__buf_1 _08328_ (.A(_04432_),
    .X(_04445_));
 sky130_fd_sc_hd__clkbuf_2 _08329_ (.A(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_1 _08330_ (.A(_04446_),
    .X(_02303_));
 sky130_fd_sc_hd__a22o_1 _08331_ (.A1(\r1.regblock[13][3] ),
    .A2(_04443_),
    .B1(_04328_),
    .B2(_04444_),
    .X(_03328_));
 sky130_fd_sc_hd__clkbuf_1 _08332_ (.A(_04446_),
    .X(_02302_));
 sky130_fd_sc_hd__a22o_1 _08333_ (.A1(\r1.regblock[13][2] ),
    .A2(_04443_),
    .B1(_04333_),
    .B2(_04444_),
    .X(_03327_));
 sky130_fd_sc_hd__clkbuf_1 _08334_ (.A(_04446_),
    .X(_02301_));
 sky130_fd_sc_hd__a22o_1 _08335_ (.A1(\r1.regblock[13][1] ),
    .A2(_04398_),
    .B1(_04335_),
    .B2(_04401_),
    .X(_03326_));
 sky130_fd_sc_hd__buf_1 _08336_ (.A(_04445_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_1 _08337_ (.A(_04447_),
    .X(_02300_));
 sky130_fd_sc_hd__a22o_1 _08338_ (.A1(\r1.regblock[13][0] ),
    .A2(_04398_),
    .B1(_04337_),
    .B2(_04401_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_1 _08339_ (.A(_04447_),
    .X(_02299_));
 sky130_fd_sc_hd__or3_1 _08340_ (.A(\r1.waddr[0] ),
    .B(_04218_),
    .C(_04221_),
    .X(_04448_));
 sky130_fd_sc_hd__buf_1 _08341_ (.A(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__or2_2 _08342_ (.A(_04394_),
    .B(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__buf_1 _08343_ (.A(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__buf_1 _08344_ (.A(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__buf_1 _08345_ (.A(\r1.wdata[31] ),
    .X(_04453_));
 sky130_fd_sc_hd__buf_1 _08346_ (.A(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__buf_1 _08347_ (.A(_04454_),
    .X(_04455_));
 sky130_fd_sc_hd__inv_2 _08348_ (.A(_04450_),
    .Y(_04456_));
 sky130_fd_sc_hd__buf_1 _08349_ (.A(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__buf_1 _08350_ (.A(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__a22o_1 _08351_ (.A1(\r1.regblock[14][31] ),
    .A2(_04452_),
    .B1(_04455_),
    .B2(_04458_),
    .X(_03324_));
 sky130_fd_sc_hd__clkbuf_1 _08352_ (.A(_04447_),
    .X(_02298_));
 sky130_fd_sc_hd__buf_1 _08353_ (.A(\r1.wdata[30] ),
    .X(_04459_));
 sky130_fd_sc_hd__buf_1 _08354_ (.A(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__buf_1 _08355_ (.A(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__a22o_1 _08356_ (.A1(\r1.regblock[14][30] ),
    .A2(_04452_),
    .B1(_04461_),
    .B2(_04458_),
    .X(_03323_));
 sky130_fd_sc_hd__buf_2 _08357_ (.A(_04445_),
    .X(_04462_));
 sky130_fd_sc_hd__clkbuf_1 _08358_ (.A(_04462_),
    .X(_02297_));
 sky130_fd_sc_hd__buf_1 _08359_ (.A(\r1.wdata[29] ),
    .X(_04463_));
 sky130_fd_sc_hd__buf_1 _08360_ (.A(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__buf_1 _08361_ (.A(_04464_),
    .X(_04465_));
 sky130_fd_sc_hd__a22o_1 _08362_ (.A1(\r1.regblock[14][29] ),
    .A2(_04452_),
    .B1(_04465_),
    .B2(_04458_),
    .X(_03322_));
 sky130_fd_sc_hd__clkbuf_1 _08363_ (.A(_04462_),
    .X(_02296_));
 sky130_fd_sc_hd__buf_4 _08364_ (.A(_04450_),
    .X(_04466_));
 sky130_fd_sc_hd__clkbuf_2 _08365_ (.A(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__buf_1 _08366_ (.A(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__buf_1 _08367_ (.A(\r1.wdata[28] ),
    .X(_04469_));
 sky130_fd_sc_hd__buf_1 _08368_ (.A(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__buf_1 _08369_ (.A(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__buf_4 _08370_ (.A(_04456_),
    .X(_04472_));
 sky130_fd_sc_hd__clkbuf_2 _08371_ (.A(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__buf_1 _08372_ (.A(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__a22o_1 _08373_ (.A1(\r1.regblock[14][28] ),
    .A2(_04468_),
    .B1(_04471_),
    .B2(_04474_),
    .X(_03321_));
 sky130_fd_sc_hd__clkbuf_1 _08374_ (.A(_04462_),
    .X(_02295_));
 sky130_fd_sc_hd__buf_1 _08375_ (.A(\r1.wdata[27] ),
    .X(_04475_));
 sky130_fd_sc_hd__clkbuf_2 _08376_ (.A(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__buf_1 _08377_ (.A(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__a22o_1 _08378_ (.A1(\r1.regblock[14][27] ),
    .A2(_04468_),
    .B1(_04477_),
    .B2(_04474_),
    .X(_03320_));
 sky130_fd_sc_hd__buf_1 _08379_ (.A(_04432_),
    .X(_04478_));
 sky130_fd_sc_hd__clkbuf_2 _08380_ (.A(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _08381_ (.A(_04479_),
    .X(_02294_));
 sky130_fd_sc_hd__buf_1 _08382_ (.A(\r1.wdata[26] ),
    .X(_04480_));
 sky130_fd_sc_hd__clkbuf_2 _08383_ (.A(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__buf_1 _08384_ (.A(_04481_),
    .X(_04482_));
 sky130_fd_sc_hd__a22o_1 _08385_ (.A1(\r1.regblock[14][26] ),
    .A2(_04468_),
    .B1(_04482_),
    .B2(_04474_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_1 _08386_ (.A(_04479_),
    .X(_02293_));
 sky130_fd_sc_hd__buf_1 _08387_ (.A(_04467_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_2 _08388_ (.A(\r1.wdata[25] ),
    .X(_04484_));
 sky130_fd_sc_hd__buf_1 _08389_ (.A(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__buf_1 _08390_ (.A(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__buf_1 _08391_ (.A(_04473_),
    .X(_04487_));
 sky130_fd_sc_hd__a22o_1 _08392_ (.A1(\r1.regblock[14][25] ),
    .A2(_04483_),
    .B1(_04486_),
    .B2(_04487_),
    .X(_03318_));
 sky130_fd_sc_hd__clkbuf_1 _08393_ (.A(_04479_),
    .X(_02292_));
 sky130_fd_sc_hd__buf_1 _08394_ (.A(\r1.wdata[24] ),
    .X(_04488_));
 sky130_fd_sc_hd__buf_1 _08395_ (.A(_04488_),
    .X(_04489_));
 sky130_fd_sc_hd__buf_1 _08396_ (.A(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__a22o_1 _08397_ (.A1(\r1.regblock[14][24] ),
    .A2(_04483_),
    .B1(_04490_),
    .B2(_04487_),
    .X(_03317_));
 sky130_fd_sc_hd__buf_1 _08398_ (.A(_04478_),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _08399_ (.A(_04491_),
    .X(_02291_));
 sky130_fd_sc_hd__clkbuf_2 _08400_ (.A(\r1.wdata[23] ),
    .X(_04492_));
 sky130_fd_sc_hd__buf_1 _08401_ (.A(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__buf_1 _08402_ (.A(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__a22o_1 _08403_ (.A1(\r1.regblock[14][23] ),
    .A2(_04483_),
    .B1(_04494_),
    .B2(_04487_),
    .X(_03316_));
 sky130_fd_sc_hd__clkbuf_1 _08404_ (.A(_04491_),
    .X(_02290_));
 sky130_fd_sc_hd__buf_1 _08405_ (.A(_04467_),
    .X(_04495_));
 sky130_fd_sc_hd__buf_1 _08406_ (.A(\r1.wdata[22] ),
    .X(_04496_));
 sky130_fd_sc_hd__buf_1 _08407_ (.A(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__buf_1 _08408_ (.A(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__buf_1 _08409_ (.A(_04473_),
    .X(_04499_));
 sky130_fd_sc_hd__a22o_1 _08410_ (.A1(\r1.regblock[14][22] ),
    .A2(_04495_),
    .B1(_04498_),
    .B2(_04499_),
    .X(_03315_));
 sky130_fd_sc_hd__clkbuf_1 _08411_ (.A(_04491_),
    .X(_02289_));
 sky130_fd_sc_hd__buf_1 _08412_ (.A(\r1.wdata[21] ),
    .X(_04500_));
 sky130_fd_sc_hd__buf_1 _08413_ (.A(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__buf_1 _08414_ (.A(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__a22o_1 _08415_ (.A1(\r1.regblock[14][21] ),
    .A2(_04495_),
    .B1(_04502_),
    .B2(_04499_),
    .X(_03314_));
 sky130_fd_sc_hd__clkbuf_4 _08416_ (.A(_04478_),
    .X(_04503_));
 sky130_fd_sc_hd__clkbuf_1 _08417_ (.A(_04503_),
    .X(_02288_));
 sky130_fd_sc_hd__buf_1 _08418_ (.A(\r1.wdata[20] ),
    .X(_04504_));
 sky130_fd_sc_hd__buf_1 _08419_ (.A(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__buf_1 _08420_ (.A(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__a22o_1 _08421_ (.A1(\r1.regblock[14][20] ),
    .A2(_04495_),
    .B1(_04506_),
    .B2(_04499_),
    .X(_03313_));
 sky130_fd_sc_hd__clkbuf_1 _08422_ (.A(_04503_),
    .X(_02287_));
 sky130_fd_sc_hd__clkbuf_2 _08423_ (.A(_04466_),
    .X(_04507_));
 sky130_fd_sc_hd__buf_1 _08424_ (.A(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__buf_1 _08425_ (.A(\r1.wdata[19] ),
    .X(_04509_));
 sky130_fd_sc_hd__buf_1 _08426_ (.A(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__buf_1 _08427_ (.A(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__clkbuf_2 _08428_ (.A(_04472_),
    .X(_04512_));
 sky130_fd_sc_hd__buf_1 _08429_ (.A(_04512_),
    .X(_04513_));
 sky130_fd_sc_hd__a22o_1 _08430_ (.A1(\r1.regblock[14][19] ),
    .A2(_04508_),
    .B1(_04511_),
    .B2(_04513_),
    .X(_03312_));
 sky130_fd_sc_hd__clkbuf_1 _08431_ (.A(_04503_),
    .X(_02286_));
 sky130_fd_sc_hd__buf_1 _08432_ (.A(\r1.wdata[18] ),
    .X(_04514_));
 sky130_fd_sc_hd__buf_1 _08433_ (.A(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__buf_1 _08434_ (.A(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__a22o_1 _08435_ (.A1(\r1.regblock[14][18] ),
    .A2(_04508_),
    .B1(_04516_),
    .B2(_04513_),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_2 _08436_ (.A(_04431_),
    .X(_04517_));
 sky130_fd_sc_hd__clkbuf_4 _08437_ (.A(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__buf_1 _08438_ (.A(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _08439_ (.A(_04519_),
    .X(_02285_));
 sky130_fd_sc_hd__buf_1 _08440_ (.A(\r1.wdata[17] ),
    .X(_04520_));
 sky130_fd_sc_hd__buf_1 _08441_ (.A(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__buf_1 _08442_ (.A(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__a22o_1 _08443_ (.A1(\r1.regblock[14][17] ),
    .A2(_04508_),
    .B1(_04522_),
    .B2(_04513_),
    .X(_03310_));
 sky130_fd_sc_hd__clkbuf_1 _08444_ (.A(_04519_),
    .X(_02284_));
 sky130_fd_sc_hd__buf_1 _08445_ (.A(_04507_),
    .X(_04523_));
 sky130_fd_sc_hd__buf_1 _08446_ (.A(\r1.wdata[16] ),
    .X(_04524_));
 sky130_fd_sc_hd__buf_1 _08447_ (.A(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__buf_1 _08448_ (.A(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__buf_1 _08449_ (.A(_04512_),
    .X(_04527_));
 sky130_fd_sc_hd__a22o_1 _08450_ (.A1(\r1.regblock[14][16] ),
    .A2(_04523_),
    .B1(_04526_),
    .B2(_04527_),
    .X(_03309_));
 sky130_fd_sc_hd__clkbuf_1 _08451_ (.A(_04519_),
    .X(_02283_));
 sky130_fd_sc_hd__buf_1 _08452_ (.A(\r1.wdata[15] ),
    .X(_04528_));
 sky130_fd_sc_hd__buf_1 _08453_ (.A(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__buf_1 _08454_ (.A(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__a22o_1 _08455_ (.A1(\r1.regblock[14][15] ),
    .A2(_04523_),
    .B1(_04530_),
    .B2(_04527_),
    .X(_03308_));
 sky130_fd_sc_hd__buf_1 _08456_ (.A(_04518_),
    .X(_04531_));
 sky130_fd_sc_hd__clkbuf_1 _08457_ (.A(_04531_),
    .X(_02282_));
 sky130_fd_sc_hd__buf_1 _08458_ (.A(\r1.wdata[14] ),
    .X(_04532_));
 sky130_fd_sc_hd__clkbuf_2 _08459_ (.A(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__buf_1 _08460_ (.A(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__a22o_1 _08461_ (.A1(\r1.regblock[14][14] ),
    .A2(_04523_),
    .B1(_04534_),
    .B2(_04527_),
    .X(_03307_));
 sky130_fd_sc_hd__clkbuf_1 _08462_ (.A(_04531_),
    .X(_02281_));
 sky130_fd_sc_hd__buf_1 _08463_ (.A(_04507_),
    .X(_04535_));
 sky130_fd_sc_hd__buf_1 _08464_ (.A(\r1.wdata[13] ),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_2 _08465_ (.A(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__buf_1 _08466_ (.A(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__buf_1 _08467_ (.A(_04512_),
    .X(_04539_));
 sky130_fd_sc_hd__a22o_1 _08468_ (.A1(\r1.regblock[14][13] ),
    .A2(_04535_),
    .B1(_04538_),
    .B2(_04539_),
    .X(_03306_));
 sky130_fd_sc_hd__clkbuf_1 _08469_ (.A(_04531_),
    .X(_02280_));
 sky130_fd_sc_hd__buf_1 _08470_ (.A(\r1.wdata[12] ),
    .X(_04540_));
 sky130_fd_sc_hd__clkbuf_2 _08471_ (.A(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__buf_1 _08472_ (.A(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__a22o_1 _08473_ (.A1(\r1.regblock[14][12] ),
    .A2(_04535_),
    .B1(_04542_),
    .B2(_04539_),
    .X(_03305_));
 sky130_fd_sc_hd__buf_2 _08474_ (.A(_04518_),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_1 _08475_ (.A(_04543_),
    .X(_02279_));
 sky130_fd_sc_hd__buf_1 _08476_ (.A(\r1.wdata[11] ),
    .X(_04544_));
 sky130_fd_sc_hd__buf_1 _08477_ (.A(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__buf_1 _08478_ (.A(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__a22o_1 _08479_ (.A1(\r1.regblock[14][11] ),
    .A2(_04535_),
    .B1(_04546_),
    .B2(_04539_),
    .X(_03304_));
 sky130_fd_sc_hd__clkbuf_1 _08480_ (.A(_04543_),
    .X(_02278_));
 sky130_fd_sc_hd__buf_1 _08481_ (.A(_04466_),
    .X(_04547_));
 sky130_fd_sc_hd__buf_1 _08482_ (.A(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__buf_1 _08483_ (.A(\r1.wdata[10] ),
    .X(_04549_));
 sky130_fd_sc_hd__buf_1 _08484_ (.A(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__buf_1 _08485_ (.A(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__buf_1 _08486_ (.A(_04472_),
    .X(_04552_));
 sky130_fd_sc_hd__buf_1 _08487_ (.A(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__a22o_1 _08488_ (.A1(\r1.regblock[14][10] ),
    .A2(_04548_),
    .B1(_04551_),
    .B2(_04553_),
    .X(_03303_));
 sky130_fd_sc_hd__clkbuf_1 _08489_ (.A(_04543_),
    .X(_02277_));
 sky130_fd_sc_hd__buf_1 _08490_ (.A(\r1.wdata[9] ),
    .X(_04554_));
 sky130_fd_sc_hd__buf_1 _08491_ (.A(_04554_),
    .X(_04555_));
 sky130_fd_sc_hd__buf_1 _08492_ (.A(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__a22o_1 _08493_ (.A1(\r1.regblock[14][9] ),
    .A2(_04548_),
    .B1(_04556_),
    .B2(_04553_),
    .X(_03302_));
 sky130_fd_sc_hd__buf_1 _08494_ (.A(_04517_),
    .X(_04557_));
 sky130_fd_sc_hd__buf_1 _08495_ (.A(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__clkbuf_1 _08496_ (.A(_04558_),
    .X(_02276_));
 sky130_fd_sc_hd__buf_1 _08497_ (.A(\r1.wdata[8] ),
    .X(_04559_));
 sky130_fd_sc_hd__buf_1 _08498_ (.A(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__buf_1 _08499_ (.A(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__a22o_1 _08500_ (.A1(\r1.regblock[14][8] ),
    .A2(_04548_),
    .B1(_04561_),
    .B2(_04553_),
    .X(_03301_));
 sky130_fd_sc_hd__clkbuf_1 _08501_ (.A(_04558_),
    .X(_02275_));
 sky130_fd_sc_hd__buf_1 _08502_ (.A(_04547_),
    .X(_04562_));
 sky130_fd_sc_hd__buf_1 _08503_ (.A(\r1.wdata[7] ),
    .X(_04563_));
 sky130_fd_sc_hd__buf_1 _08504_ (.A(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__buf_1 _08505_ (.A(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__buf_1 _08506_ (.A(_04552_),
    .X(_04566_));
 sky130_fd_sc_hd__a22o_1 _08507_ (.A1(\r1.regblock[14][7] ),
    .A2(_04562_),
    .B1(_04565_),
    .B2(_04566_),
    .X(_03300_));
 sky130_fd_sc_hd__clkbuf_1 _08508_ (.A(_04558_),
    .X(_02274_));
 sky130_fd_sc_hd__buf_1 _08509_ (.A(\r1.wdata[6] ),
    .X(_04567_));
 sky130_fd_sc_hd__buf_1 _08510_ (.A(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__buf_1 _08511_ (.A(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__a22o_1 _08512_ (.A1(\r1.regblock[14][6] ),
    .A2(_04562_),
    .B1(_04569_),
    .B2(_04566_),
    .X(_03299_));
 sky130_fd_sc_hd__buf_1 _08513_ (.A(_04557_),
    .X(_04570_));
 sky130_fd_sc_hd__clkbuf_1 _08514_ (.A(_04570_),
    .X(_02273_));
 sky130_fd_sc_hd__buf_1 _08515_ (.A(\r1.wdata[5] ),
    .X(_04571_));
 sky130_fd_sc_hd__buf_1 _08516_ (.A(_04571_),
    .X(_04572_));
 sky130_fd_sc_hd__buf_1 _08517_ (.A(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__a22o_1 _08518_ (.A1(\r1.regblock[14][5] ),
    .A2(_04562_),
    .B1(_04573_),
    .B2(_04566_),
    .X(_03298_));
 sky130_fd_sc_hd__clkbuf_1 _08519_ (.A(_04570_),
    .X(_02272_));
 sky130_fd_sc_hd__buf_1 _08520_ (.A(_04547_),
    .X(_04574_));
 sky130_fd_sc_hd__buf_1 _08521_ (.A(\r1.wdata[4] ),
    .X(_04575_));
 sky130_fd_sc_hd__buf_1 _08522_ (.A(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__buf_1 _08523_ (.A(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__buf_1 _08524_ (.A(_04552_),
    .X(_04578_));
 sky130_fd_sc_hd__a22o_1 _08525_ (.A1(\r1.regblock[14][4] ),
    .A2(_04574_),
    .B1(_04577_),
    .B2(_04578_),
    .X(_03297_));
 sky130_fd_sc_hd__clkbuf_1 _08526_ (.A(_04570_),
    .X(_02271_));
 sky130_fd_sc_hd__buf_1 _08527_ (.A(\r1.wdata[3] ),
    .X(_04579_));
 sky130_fd_sc_hd__buf_1 _08528_ (.A(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__buf_1 _08529_ (.A(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__a22o_1 _08530_ (.A1(\r1.regblock[14][3] ),
    .A2(_04574_),
    .B1(_04581_),
    .B2(_04578_),
    .X(_03296_));
 sky130_fd_sc_hd__buf_2 _08531_ (.A(_04557_),
    .X(_04582_));
 sky130_fd_sc_hd__clkbuf_1 _08532_ (.A(_04582_),
    .X(_02270_));
 sky130_fd_sc_hd__buf_1 _08533_ (.A(\r1.wdata[2] ),
    .X(_04583_));
 sky130_fd_sc_hd__clkbuf_2 _08534_ (.A(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__buf_1 _08535_ (.A(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__a22o_1 _08536_ (.A1(\r1.regblock[14][2] ),
    .A2(_04574_),
    .B1(_04585_),
    .B2(_04578_),
    .X(_03295_));
 sky130_fd_sc_hd__clkbuf_1 _08537_ (.A(_04582_),
    .X(_02269_));
 sky130_fd_sc_hd__buf_1 _08538_ (.A(\r1.wdata[1] ),
    .X(_04586_));
 sky130_fd_sc_hd__buf_1 _08539_ (.A(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__buf_1 _08540_ (.A(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__a22o_1 _08541_ (.A1(\r1.regblock[14][1] ),
    .A2(_04451_),
    .B1(_04588_),
    .B2(_04457_),
    .X(_03294_));
 sky130_fd_sc_hd__clkbuf_1 _08542_ (.A(_04582_),
    .X(_02268_));
 sky130_fd_sc_hd__buf_1 _08543_ (.A(\r1.wdata[0] ),
    .X(_04589_));
 sky130_fd_sc_hd__buf_1 _08544_ (.A(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__buf_1 _08545_ (.A(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__a22o_1 _08546_ (.A1(\r1.regblock[14][0] ),
    .A2(_04451_),
    .B1(_04591_),
    .B2(_04457_),
    .X(_03293_));
 sky130_fd_sc_hd__clkbuf_4 _08547_ (.A(_04517_),
    .X(_04592_));
 sky130_fd_sc_hd__buf_1 _08548_ (.A(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__clkbuf_1 _08549_ (.A(_04593_),
    .X(_02267_));
 sky130_fd_sc_hd__or2_2 _08550_ (.A(_04339_),
    .B(_04393_),
    .X(_04594_));
 sky130_fd_sc_hd__buf_1 _08551_ (.A(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__buf_1 _08552_ (.A(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__inv_2 _08553_ (.A(_04594_),
    .Y(_04597_));
 sky130_fd_sc_hd__buf_1 _08554_ (.A(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__buf_1 _08555_ (.A(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__a22o_1 _08556_ (.A1(\r1.regblock[15][31] ),
    .A2(_04596_),
    .B1(_04455_),
    .B2(_04599_),
    .X(_03292_));
 sky130_fd_sc_hd__clkbuf_1 _08557_ (.A(_04593_),
    .X(_02266_));
 sky130_fd_sc_hd__a22o_1 _08558_ (.A1(\r1.regblock[15][30] ),
    .A2(_04596_),
    .B1(_04461_),
    .B2(_04599_),
    .X(_03291_));
 sky130_fd_sc_hd__clkbuf_1 _08559_ (.A(_04593_),
    .X(_02265_));
 sky130_fd_sc_hd__a22o_1 _08560_ (.A1(\r1.regblock[15][29] ),
    .A2(_04596_),
    .B1(_04465_),
    .B2(_04599_),
    .X(_03290_));
 sky130_fd_sc_hd__buf_1 _08561_ (.A(_04592_),
    .X(_04600_));
 sky130_fd_sc_hd__clkbuf_1 _08562_ (.A(_04600_),
    .X(_02264_));
 sky130_fd_sc_hd__clkbuf_4 _08563_ (.A(_04594_),
    .X(_04601_));
 sky130_fd_sc_hd__clkbuf_2 _08564_ (.A(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__buf_1 _08565_ (.A(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__clkbuf_4 _08566_ (.A(_04597_),
    .X(_04604_));
 sky130_fd_sc_hd__clkbuf_2 _08567_ (.A(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__buf_1 _08568_ (.A(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__a22o_1 _08569_ (.A1(\r1.regblock[15][28] ),
    .A2(_04603_),
    .B1(_04471_),
    .B2(_04606_),
    .X(_03289_));
 sky130_fd_sc_hd__clkbuf_1 _08570_ (.A(_04600_),
    .X(_02263_));
 sky130_fd_sc_hd__a22o_1 _08571_ (.A1(\r1.regblock[15][27] ),
    .A2(_04603_),
    .B1(_04477_),
    .B2(_04606_),
    .X(_03288_));
 sky130_fd_sc_hd__clkbuf_1 _08572_ (.A(_04600_),
    .X(_02262_));
 sky130_fd_sc_hd__a22o_1 _08573_ (.A1(\r1.regblock[15][26] ),
    .A2(_04603_),
    .B1(_04482_),
    .B2(_04606_),
    .X(_03287_));
 sky130_fd_sc_hd__buf_1 _08574_ (.A(_04592_),
    .X(_04607_));
 sky130_fd_sc_hd__clkbuf_1 _08575_ (.A(_04607_),
    .X(_02261_));
 sky130_fd_sc_hd__buf_1 _08576_ (.A(_04602_),
    .X(_04608_));
 sky130_fd_sc_hd__buf_1 _08577_ (.A(_04605_),
    .X(_04609_));
 sky130_fd_sc_hd__a22o_1 _08578_ (.A1(\r1.regblock[15][25] ),
    .A2(_04608_),
    .B1(_04486_),
    .B2(_04609_),
    .X(_03286_));
 sky130_fd_sc_hd__clkbuf_1 _08579_ (.A(_04607_),
    .X(_02260_));
 sky130_fd_sc_hd__a22o_1 _08580_ (.A1(\r1.regblock[15][24] ),
    .A2(_04608_),
    .B1(_04490_),
    .B2(_04609_),
    .X(_03285_));
 sky130_fd_sc_hd__clkbuf_1 _08581_ (.A(_04607_),
    .X(_02259_));
 sky130_fd_sc_hd__a22o_1 _08582_ (.A1(\r1.regblock[15][23] ),
    .A2(_04608_),
    .B1(_04494_),
    .B2(_04609_),
    .X(_03284_));
 sky130_fd_sc_hd__buf_1 _08583_ (.A(_04431_),
    .X(_04610_));
 sky130_fd_sc_hd__clkbuf_4 _08584_ (.A(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__buf_1 _08585_ (.A(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__clkbuf_1 _08586_ (.A(_04612_),
    .X(_02258_));
 sky130_fd_sc_hd__buf_1 _08587_ (.A(_04602_),
    .X(_04613_));
 sky130_fd_sc_hd__buf_1 _08588_ (.A(_04605_),
    .X(_04614_));
 sky130_fd_sc_hd__a22o_1 _08589_ (.A1(\r1.regblock[15][22] ),
    .A2(_04613_),
    .B1(_04498_),
    .B2(_04614_),
    .X(_03283_));
 sky130_fd_sc_hd__clkbuf_1 _08590_ (.A(_04612_),
    .X(_02257_));
 sky130_fd_sc_hd__a22o_1 _08591_ (.A1(\r1.regblock[15][21] ),
    .A2(_04613_),
    .B1(_04502_),
    .B2(_04614_),
    .X(_03282_));
 sky130_fd_sc_hd__clkbuf_1 _08592_ (.A(_04612_),
    .X(_02256_));
 sky130_fd_sc_hd__a22o_1 _08593_ (.A1(\r1.regblock[15][20] ),
    .A2(_04613_),
    .B1(_04506_),
    .B2(_04614_),
    .X(_03281_));
 sky130_fd_sc_hd__buf_1 _08594_ (.A(_04611_),
    .X(_04615_));
 sky130_fd_sc_hd__clkbuf_1 _08595_ (.A(_04615_),
    .X(_02255_));
 sky130_fd_sc_hd__clkbuf_2 _08596_ (.A(_04601_),
    .X(_04616_));
 sky130_fd_sc_hd__buf_1 _08597_ (.A(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__clkbuf_2 _08598_ (.A(_04604_),
    .X(_04618_));
 sky130_fd_sc_hd__buf_1 _08599_ (.A(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__a22o_1 _08600_ (.A1(\r1.regblock[15][19] ),
    .A2(_04617_),
    .B1(_04511_),
    .B2(_04619_),
    .X(_03280_));
 sky130_fd_sc_hd__clkbuf_1 _08601_ (.A(_04615_),
    .X(_02254_));
 sky130_fd_sc_hd__a22o_1 _08602_ (.A1(\r1.regblock[15][18] ),
    .A2(_04617_),
    .B1(_04516_),
    .B2(_04619_),
    .X(_03279_));
 sky130_fd_sc_hd__clkbuf_1 _08603_ (.A(_04615_),
    .X(_02253_));
 sky130_fd_sc_hd__a22o_1 _08604_ (.A1(\r1.regblock[15][17] ),
    .A2(_04617_),
    .B1(_04522_),
    .B2(_04619_),
    .X(_03278_));
 sky130_fd_sc_hd__buf_1 _08605_ (.A(_04611_),
    .X(_04620_));
 sky130_fd_sc_hd__clkbuf_1 _08606_ (.A(_04620_),
    .X(_02252_));
 sky130_fd_sc_hd__buf_1 _08607_ (.A(_04616_),
    .X(_04621_));
 sky130_fd_sc_hd__buf_1 _08608_ (.A(_04618_),
    .X(_04622_));
 sky130_fd_sc_hd__a22o_1 _08609_ (.A1(\r1.regblock[15][16] ),
    .A2(_04621_),
    .B1(_04526_),
    .B2(_04622_),
    .X(_03277_));
 sky130_fd_sc_hd__clkbuf_1 _08610_ (.A(_04620_),
    .X(_02251_));
 sky130_fd_sc_hd__a22o_1 _08611_ (.A1(\r1.regblock[15][15] ),
    .A2(_04621_),
    .B1(_04530_),
    .B2(_04622_),
    .X(_03276_));
 sky130_fd_sc_hd__clkbuf_1 _08612_ (.A(_04620_),
    .X(_02250_));
 sky130_fd_sc_hd__a22o_1 _08613_ (.A1(\r1.regblock[15][14] ),
    .A2(_04621_),
    .B1(_04534_),
    .B2(_04622_),
    .X(_03275_));
 sky130_fd_sc_hd__buf_4 _08614_ (.A(_04610_),
    .X(_04623_));
 sky130_fd_sc_hd__buf_1 _08615_ (.A(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__clkbuf_1 _08616_ (.A(_04624_),
    .X(_02249_));
 sky130_fd_sc_hd__buf_1 _08617_ (.A(_04616_),
    .X(_04625_));
 sky130_fd_sc_hd__buf_1 _08618_ (.A(_04618_),
    .X(_04626_));
 sky130_fd_sc_hd__a22o_1 _08619_ (.A1(\r1.regblock[15][13] ),
    .A2(_04625_),
    .B1(_04538_),
    .B2(_04626_),
    .X(_03274_));
 sky130_fd_sc_hd__clkbuf_1 _08620_ (.A(_04624_),
    .X(_02248_));
 sky130_fd_sc_hd__a22o_1 _08621_ (.A1(\r1.regblock[15][12] ),
    .A2(_04625_),
    .B1(_04542_),
    .B2(_04626_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_1 _08622_ (.A(_04624_),
    .X(_02247_));
 sky130_fd_sc_hd__a22o_1 _08623_ (.A1(\r1.regblock[15][11] ),
    .A2(_04625_),
    .B1(_04546_),
    .B2(_04626_),
    .X(_03272_));
 sky130_fd_sc_hd__buf_1 _08624_ (.A(_04623_),
    .X(_04627_));
 sky130_fd_sc_hd__clkbuf_1 _08625_ (.A(_04627_),
    .X(_02246_));
 sky130_fd_sc_hd__buf_1 _08626_ (.A(_04601_),
    .X(_04628_));
 sky130_fd_sc_hd__buf_1 _08627_ (.A(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__buf_1 _08628_ (.A(_04604_),
    .X(_04630_));
 sky130_fd_sc_hd__buf_1 _08629_ (.A(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__a22o_1 _08630_ (.A1(\r1.regblock[15][10] ),
    .A2(_04629_),
    .B1(_04551_),
    .B2(_04631_),
    .X(_03271_));
 sky130_fd_sc_hd__clkbuf_1 _08631_ (.A(_04627_),
    .X(_02245_));
 sky130_fd_sc_hd__a22o_1 _08632_ (.A1(\r1.regblock[15][9] ),
    .A2(_04629_),
    .B1(_04556_),
    .B2(_04631_),
    .X(_03270_));
 sky130_fd_sc_hd__clkbuf_1 _08633_ (.A(_04627_),
    .X(_02244_));
 sky130_fd_sc_hd__a22o_1 _08634_ (.A1(\r1.regblock[15][8] ),
    .A2(_04629_),
    .B1(_04561_),
    .B2(_04631_),
    .X(_03269_));
 sky130_fd_sc_hd__buf_1 _08635_ (.A(_04623_),
    .X(_04632_));
 sky130_fd_sc_hd__clkbuf_1 _08636_ (.A(_04632_),
    .X(_02243_));
 sky130_fd_sc_hd__buf_1 _08637_ (.A(_04628_),
    .X(_04633_));
 sky130_fd_sc_hd__buf_1 _08638_ (.A(_04630_),
    .X(_04634_));
 sky130_fd_sc_hd__a22o_1 _08639_ (.A1(\r1.regblock[15][7] ),
    .A2(_04633_),
    .B1(_04565_),
    .B2(_04634_),
    .X(_03268_));
 sky130_fd_sc_hd__clkbuf_1 _08640_ (.A(_04632_),
    .X(_02242_));
 sky130_fd_sc_hd__a22o_1 _08641_ (.A1(\r1.regblock[15][6] ),
    .A2(_04633_),
    .B1(_04569_),
    .B2(_04634_),
    .X(_03267_));
 sky130_fd_sc_hd__clkbuf_1 _08642_ (.A(_04632_),
    .X(_02241_));
 sky130_fd_sc_hd__a22o_1 _08643_ (.A1(\r1.regblock[15][5] ),
    .A2(_04633_),
    .B1(_04573_),
    .B2(_04634_),
    .X(_03266_));
 sky130_fd_sc_hd__buf_2 _08644_ (.A(_04610_),
    .X(_04635_));
 sky130_fd_sc_hd__buf_1 _08645_ (.A(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__clkbuf_1 _08646_ (.A(_04636_),
    .X(_02240_));
 sky130_fd_sc_hd__buf_1 _08647_ (.A(_04628_),
    .X(_04637_));
 sky130_fd_sc_hd__buf_1 _08648_ (.A(_04630_),
    .X(_04638_));
 sky130_fd_sc_hd__a22o_1 _08649_ (.A1(\r1.regblock[15][4] ),
    .A2(_04637_),
    .B1(_04577_),
    .B2(_04638_),
    .X(_03265_));
 sky130_fd_sc_hd__clkbuf_1 _08650_ (.A(_04636_),
    .X(_02239_));
 sky130_fd_sc_hd__a22o_1 _08651_ (.A1(\r1.regblock[15][3] ),
    .A2(_04637_),
    .B1(_04581_),
    .B2(_04638_),
    .X(_03264_));
 sky130_fd_sc_hd__clkbuf_1 _08652_ (.A(_04636_),
    .X(_02238_));
 sky130_fd_sc_hd__a22o_1 _08653_ (.A1(\r1.regblock[15][2] ),
    .A2(_04637_),
    .B1(_04585_),
    .B2(_04638_),
    .X(_03263_));
 sky130_fd_sc_hd__buf_1 _08654_ (.A(_04635_),
    .X(_04639_));
 sky130_fd_sc_hd__clkbuf_1 _08655_ (.A(_04639_),
    .X(_02237_));
 sky130_fd_sc_hd__a22o_1 _08656_ (.A1(\r1.regblock[15][1] ),
    .A2(_04595_),
    .B1(_04588_),
    .B2(_04598_),
    .X(_03262_));
 sky130_fd_sc_hd__clkbuf_1 _08657_ (.A(_04639_),
    .X(_02236_));
 sky130_fd_sc_hd__a22o_1 _08658_ (.A1(\r1.regblock[15][0] ),
    .A2(_04595_),
    .B1(_04591_),
    .B2(_04598_),
    .X(_03261_));
 sky130_fd_sc_hd__clkbuf_1 _08659_ (.A(_04639_),
    .X(_02235_));
 sky130_fd_sc_hd__buf_1 _08660_ (.A(_04395_),
    .X(_04640_));
 sky130_fd_sc_hd__buf_1 _08661_ (.A(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__or3_1 _08662_ (.A(\r1.waddr[4] ),
    .B(\r1.waddr[3] ),
    .C(_04391_),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_1 _08663_ (.A(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__or2_2 _08664_ (.A(_04641_),
    .B(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__buf_1 _08665_ (.A(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__buf_1 _08666_ (.A(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__inv_2 _08667_ (.A(_04644_),
    .Y(_04647_));
 sky130_fd_sc_hd__buf_1 _08668_ (.A(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__buf_1 _08669_ (.A(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__a22o_1 _08670_ (.A1(\r1.regblock[5][31] ),
    .A2(_04646_),
    .B1(_04455_),
    .B2(_04649_),
    .X(_03260_));
 sky130_fd_sc_hd__buf_2 _08671_ (.A(_04635_),
    .X(_04650_));
 sky130_fd_sc_hd__clkbuf_1 _08672_ (.A(_04650_),
    .X(_02234_));
 sky130_fd_sc_hd__a22o_1 _08673_ (.A1(\r1.regblock[5][30] ),
    .A2(_04646_),
    .B1(_04461_),
    .B2(_04649_),
    .X(_03259_));
 sky130_fd_sc_hd__clkbuf_1 _08674_ (.A(_04650_),
    .X(_02233_));
 sky130_fd_sc_hd__a22o_1 _08675_ (.A1(\r1.regblock[5][29] ),
    .A2(_04646_),
    .B1(_04465_),
    .B2(_04649_),
    .X(_03258_));
 sky130_fd_sc_hd__clkbuf_1 _08676_ (.A(_04650_),
    .X(_02232_));
 sky130_fd_sc_hd__buf_4 _08677_ (.A(_04644_),
    .X(_04651_));
 sky130_fd_sc_hd__clkbuf_2 _08678_ (.A(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__buf_1 _08679_ (.A(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__buf_4 _08680_ (.A(_04647_),
    .X(_04654_));
 sky130_fd_sc_hd__clkbuf_2 _08681_ (.A(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__buf_1 _08682_ (.A(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__a22o_1 _08683_ (.A1(\r1.regblock[5][28] ),
    .A2(_04653_),
    .B1(_04471_),
    .B2(_04656_),
    .X(_03257_));
 sky130_fd_sc_hd__clkbuf_1 _08684_ (.A(_04430_),
    .X(_04657_));
 sky130_fd_sc_hd__clkbuf_4 _08685_ (.A(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__clkbuf_2 _08686_ (.A(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__clkbuf_2 _08687_ (.A(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__clkbuf_1 _08688_ (.A(_04660_),
    .X(_02231_));
 sky130_fd_sc_hd__a22o_1 _08689_ (.A1(\r1.regblock[5][27] ),
    .A2(_04653_),
    .B1(_04477_),
    .B2(_04656_),
    .X(_03256_));
 sky130_fd_sc_hd__clkbuf_1 _08690_ (.A(_04660_),
    .X(_02230_));
 sky130_fd_sc_hd__a22o_1 _08691_ (.A1(\r1.regblock[5][26] ),
    .A2(_04653_),
    .B1(_04482_),
    .B2(_04656_),
    .X(_03255_));
 sky130_fd_sc_hd__clkbuf_1 _08692_ (.A(_04660_),
    .X(_02229_));
 sky130_fd_sc_hd__buf_1 _08693_ (.A(_04652_),
    .X(_04661_));
 sky130_fd_sc_hd__buf_1 _08694_ (.A(_04655_),
    .X(_04662_));
 sky130_fd_sc_hd__a22o_1 _08695_ (.A1(\r1.regblock[5][25] ),
    .A2(_04661_),
    .B1(_04486_),
    .B2(_04662_),
    .X(_03254_));
 sky130_fd_sc_hd__buf_1 _08696_ (.A(_04659_),
    .X(_04663_));
 sky130_fd_sc_hd__clkbuf_1 _08697_ (.A(_04663_),
    .X(_02228_));
 sky130_fd_sc_hd__a22o_1 _08698_ (.A1(\r1.regblock[5][24] ),
    .A2(_04661_),
    .B1(_04490_),
    .B2(_04662_),
    .X(_03253_));
 sky130_fd_sc_hd__clkbuf_1 _08699_ (.A(_04663_),
    .X(_02227_));
 sky130_fd_sc_hd__a22o_1 _08700_ (.A1(\r1.regblock[5][23] ),
    .A2(_04661_),
    .B1(_04494_),
    .B2(_04662_),
    .X(_03252_));
 sky130_fd_sc_hd__clkbuf_1 _08701_ (.A(_04663_),
    .X(_02226_));
 sky130_fd_sc_hd__buf_1 _08702_ (.A(_04652_),
    .X(_04664_));
 sky130_fd_sc_hd__buf_1 _08703_ (.A(_04655_),
    .X(_04665_));
 sky130_fd_sc_hd__a22o_1 _08704_ (.A1(\r1.regblock[5][22] ),
    .A2(_04664_),
    .B1(_04498_),
    .B2(_04665_),
    .X(_03251_));
 sky130_fd_sc_hd__clkbuf_2 _08705_ (.A(_04659_),
    .X(_04666_));
 sky130_fd_sc_hd__clkbuf_1 _08706_ (.A(_04666_),
    .X(_02225_));
 sky130_fd_sc_hd__a22o_1 _08707_ (.A1(\r1.regblock[5][21] ),
    .A2(_04664_),
    .B1(_04502_),
    .B2(_04665_),
    .X(_03250_));
 sky130_fd_sc_hd__clkbuf_1 _08708_ (.A(_04666_),
    .X(_02224_));
 sky130_fd_sc_hd__a22o_1 _08709_ (.A1(\r1.regblock[5][20] ),
    .A2(_04664_),
    .B1(_04506_),
    .B2(_04665_),
    .X(_03249_));
 sky130_fd_sc_hd__clkbuf_2 _08710_ (.A(_04666_),
    .X(_02223_));
 sky130_fd_sc_hd__buf_1 _08711_ (.A(_04651_),
    .X(_04667_));
 sky130_fd_sc_hd__buf_1 _08712_ (.A(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__clkbuf_2 _08713_ (.A(_04654_),
    .X(_04669_));
 sky130_fd_sc_hd__buf_1 _08714_ (.A(_04669_),
    .X(_04670_));
 sky130_fd_sc_hd__a22o_1 _08715_ (.A1(\r1.regblock[5][19] ),
    .A2(_04668_),
    .B1(_04511_),
    .B2(_04670_),
    .X(_03248_));
 sky130_fd_sc_hd__buf_1 _08716_ (.A(_04658_),
    .X(_04671_));
 sky130_fd_sc_hd__buf_1 _08717_ (.A(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__clkbuf_1 _08718_ (.A(_04672_),
    .X(_02222_));
 sky130_fd_sc_hd__a22o_1 _08719_ (.A1(\r1.regblock[5][18] ),
    .A2(_04668_),
    .B1(_04516_),
    .B2(_04670_),
    .X(_03247_));
 sky130_fd_sc_hd__clkbuf_1 _08720_ (.A(_04672_),
    .X(_02221_));
 sky130_fd_sc_hd__a22o_1 _08721_ (.A1(\r1.regblock[5][17] ),
    .A2(_04668_),
    .B1(_04522_),
    .B2(_04670_),
    .X(_03246_));
 sky130_fd_sc_hd__clkbuf_1 _08722_ (.A(_04672_),
    .X(_02220_));
 sky130_fd_sc_hd__buf_1 _08723_ (.A(_04667_),
    .X(_04673_));
 sky130_fd_sc_hd__buf_1 _08724_ (.A(_04669_),
    .X(_04674_));
 sky130_fd_sc_hd__a22o_1 _08725_ (.A1(\r1.regblock[5][16] ),
    .A2(_04673_),
    .B1(_04526_),
    .B2(_04674_),
    .X(_03245_));
 sky130_fd_sc_hd__buf_1 _08726_ (.A(_04671_),
    .X(_04675_));
 sky130_fd_sc_hd__clkbuf_1 _08727_ (.A(_04675_),
    .X(_02219_));
 sky130_fd_sc_hd__a22o_1 _08728_ (.A1(\r1.regblock[5][15] ),
    .A2(_04673_),
    .B1(_04530_),
    .B2(_04674_),
    .X(_03244_));
 sky130_fd_sc_hd__clkbuf_1 _08729_ (.A(_04675_),
    .X(_02218_));
 sky130_fd_sc_hd__a22o_1 _08730_ (.A1(\r1.regblock[5][14] ),
    .A2(_04673_),
    .B1(_04534_),
    .B2(_04674_),
    .X(_03243_));
 sky130_fd_sc_hd__clkbuf_1 _08731_ (.A(_04675_),
    .X(_02217_));
 sky130_fd_sc_hd__buf_1 _08732_ (.A(_04667_),
    .X(_04676_));
 sky130_fd_sc_hd__buf_1 _08733_ (.A(_04669_),
    .X(_04677_));
 sky130_fd_sc_hd__a22o_1 _08734_ (.A1(\r1.regblock[5][13] ),
    .A2(_04676_),
    .B1(_04538_),
    .B2(_04677_),
    .X(_03242_));
 sky130_fd_sc_hd__buf_1 _08735_ (.A(_04671_),
    .X(_04678_));
 sky130_fd_sc_hd__clkbuf_1 _08736_ (.A(_04678_),
    .X(_02216_));
 sky130_fd_sc_hd__a22o_1 _08737_ (.A1(\r1.regblock[5][12] ),
    .A2(_04676_),
    .B1(_04542_),
    .B2(_04677_),
    .X(_03241_));
 sky130_fd_sc_hd__clkbuf_1 _08738_ (.A(_04678_),
    .X(_02215_));
 sky130_fd_sc_hd__a22o_1 _08739_ (.A1(\r1.regblock[5][11] ),
    .A2(_04676_),
    .B1(_04546_),
    .B2(_04677_),
    .X(_03240_));
 sky130_fd_sc_hd__clkbuf_2 _08740_ (.A(_04678_),
    .X(_02214_));
 sky130_fd_sc_hd__buf_1 _08741_ (.A(_04651_),
    .X(_04679_));
 sky130_fd_sc_hd__buf_1 _08742_ (.A(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__buf_1 _08743_ (.A(_04654_),
    .X(_04681_));
 sky130_fd_sc_hd__buf_1 _08744_ (.A(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__a22o_1 _08745_ (.A1(\r1.regblock[5][10] ),
    .A2(_04680_),
    .B1(_04551_),
    .B2(_04682_),
    .X(_03239_));
 sky130_fd_sc_hd__buf_1 _08746_ (.A(_04658_),
    .X(_04683_));
 sky130_fd_sc_hd__buf_1 _08747_ (.A(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__clkbuf_1 _08748_ (.A(_04684_),
    .X(_02213_));
 sky130_fd_sc_hd__a22o_1 _08749_ (.A1(\r1.regblock[5][9] ),
    .A2(_04680_),
    .B1(_04556_),
    .B2(_04682_),
    .X(_03238_));
 sky130_fd_sc_hd__clkbuf_1 _08750_ (.A(_04684_),
    .X(_02212_));
 sky130_fd_sc_hd__a22o_1 _08751_ (.A1(\r1.regblock[5][8] ),
    .A2(_04680_),
    .B1(_04561_),
    .B2(_04682_),
    .X(_03237_));
 sky130_fd_sc_hd__clkbuf_1 _08752_ (.A(_04684_),
    .X(_02211_));
 sky130_fd_sc_hd__buf_1 _08753_ (.A(_04679_),
    .X(_04685_));
 sky130_fd_sc_hd__buf_1 _08754_ (.A(_04681_),
    .X(_04686_));
 sky130_fd_sc_hd__a22o_1 _08755_ (.A1(\r1.regblock[5][7] ),
    .A2(_04685_),
    .B1(_04565_),
    .B2(_04686_),
    .X(_03236_));
 sky130_fd_sc_hd__buf_1 _08756_ (.A(_04683_),
    .X(_04687_));
 sky130_fd_sc_hd__clkbuf_1 _08757_ (.A(_04687_),
    .X(_02210_));
 sky130_fd_sc_hd__a22o_1 _08758_ (.A1(\r1.regblock[5][6] ),
    .A2(_04685_),
    .B1(_04569_),
    .B2(_04686_),
    .X(_03235_));
 sky130_fd_sc_hd__clkbuf_1 _08759_ (.A(_04687_),
    .X(_02209_));
 sky130_fd_sc_hd__a22o_1 _08760_ (.A1(\r1.regblock[5][5] ),
    .A2(_04685_),
    .B1(_04573_),
    .B2(_04686_),
    .X(_03234_));
 sky130_fd_sc_hd__clkbuf_1 _08761_ (.A(_04687_),
    .X(_02208_));
 sky130_fd_sc_hd__buf_1 _08762_ (.A(_04679_),
    .X(_04688_));
 sky130_fd_sc_hd__buf_1 _08763_ (.A(_04681_),
    .X(_04689_));
 sky130_fd_sc_hd__a22o_1 _08764_ (.A1(\r1.regblock[5][4] ),
    .A2(_04688_),
    .B1(_04577_),
    .B2(_04689_),
    .X(_03233_));
 sky130_fd_sc_hd__buf_1 _08765_ (.A(_04683_),
    .X(_04690_));
 sky130_fd_sc_hd__clkbuf_1 _08766_ (.A(_04690_),
    .X(_02207_));
 sky130_fd_sc_hd__a22o_1 _08767_ (.A1(\r1.regblock[5][3] ),
    .A2(_04688_),
    .B1(_04581_),
    .B2(_04689_),
    .X(_03232_));
 sky130_fd_sc_hd__clkbuf_1 _08768_ (.A(_04690_),
    .X(_02206_));
 sky130_fd_sc_hd__a22o_1 _08769_ (.A1(\r1.regblock[5][2] ),
    .A2(_04688_),
    .B1(_04585_),
    .B2(_04689_),
    .X(_03231_));
 sky130_fd_sc_hd__clkbuf_2 _08770_ (.A(_04690_),
    .X(_02205_));
 sky130_fd_sc_hd__a22o_1 _08771_ (.A1(\r1.regblock[5][1] ),
    .A2(_04645_),
    .B1(_04588_),
    .B2(_04648_),
    .X(_03230_));
 sky130_fd_sc_hd__buf_2 _08772_ (.A(_04657_),
    .X(_04691_));
 sky130_fd_sc_hd__buf_1 _08773_ (.A(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__buf_1 _08774_ (.A(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__clkbuf_1 _08775_ (.A(_04693_),
    .X(_02204_));
 sky130_fd_sc_hd__a22o_1 _08776_ (.A1(\r1.regblock[5][0] ),
    .A2(_04645_),
    .B1(_04591_),
    .B2(_04648_),
    .X(_03229_));
 sky130_fd_sc_hd__clkbuf_1 _08777_ (.A(_04693_),
    .X(_02203_));
 sky130_fd_sc_hd__or3_1 _08778_ (.A(\r1.waddr[0] ),
    .B(\r1.waddr[1] ),
    .C(_04221_),
    .X(_04694_));
 sky130_fd_sc_hd__buf_1 _08779_ (.A(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__or2_2 _08780_ (.A(_04217_),
    .B(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__buf_1 _08781_ (.A(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__buf_1 _08782_ (.A(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__buf_1 _08783_ (.A(_04454_),
    .X(_04699_));
 sky130_fd_sc_hd__inv_2 _08784_ (.A(_04696_),
    .Y(_04700_));
 sky130_fd_sc_hd__buf_1 _08785_ (.A(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__buf_1 _08786_ (.A(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__a22o_1 _08787_ (.A1(\r1.regblock[0][31] ),
    .A2(_04698_),
    .B1(_04699_),
    .B2(_04702_),
    .X(_03228_));
 sky130_fd_sc_hd__clkbuf_1 _08788_ (.A(_04693_),
    .X(_02202_));
 sky130_fd_sc_hd__buf_1 _08789_ (.A(_04460_),
    .X(_04703_));
 sky130_fd_sc_hd__a22o_1 _08790_ (.A1(\r1.regblock[0][30] ),
    .A2(_04698_),
    .B1(_04703_),
    .B2(_04702_),
    .X(_03227_));
 sky130_fd_sc_hd__clkbuf_2 _08791_ (.A(_04692_),
    .X(_04704_));
 sky130_fd_sc_hd__clkbuf_1 _08792_ (.A(_04704_),
    .X(_02201_));
 sky130_fd_sc_hd__buf_1 _08793_ (.A(_04464_),
    .X(_04705_));
 sky130_fd_sc_hd__a22o_1 _08794_ (.A1(\r1.regblock[0][29] ),
    .A2(_04698_),
    .B1(_04705_),
    .B2(_04702_),
    .X(_03226_));
 sky130_fd_sc_hd__clkbuf_1 _08795_ (.A(_04704_),
    .X(_02200_));
 sky130_fd_sc_hd__clkbuf_4 _08796_ (.A(_04696_),
    .X(_04706_));
 sky130_fd_sc_hd__clkbuf_2 _08797_ (.A(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__buf_1 _08798_ (.A(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__buf_1 _08799_ (.A(_04470_),
    .X(_04709_));
 sky130_fd_sc_hd__clkbuf_4 _08800_ (.A(_04700_),
    .X(_04710_));
 sky130_fd_sc_hd__clkbuf_2 _08801_ (.A(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__buf_1 _08802_ (.A(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__a22o_1 _08803_ (.A1(\r1.regblock[0][28] ),
    .A2(_04708_),
    .B1(_04709_),
    .B2(_04712_),
    .X(_03225_));
 sky130_fd_sc_hd__clkbuf_1 _08804_ (.A(_04704_),
    .X(_02199_));
 sky130_fd_sc_hd__buf_1 _08805_ (.A(_04476_),
    .X(_04713_));
 sky130_fd_sc_hd__a22o_1 _08806_ (.A1(\r1.regblock[0][27] ),
    .A2(_04708_),
    .B1(_04713_),
    .B2(_04712_),
    .X(_03224_));
 sky130_fd_sc_hd__buf_1 _08807_ (.A(_04692_),
    .X(_04714_));
 sky130_fd_sc_hd__clkbuf_1 _08808_ (.A(_04714_),
    .X(_02198_));
 sky130_fd_sc_hd__buf_1 _08809_ (.A(_04481_),
    .X(_04715_));
 sky130_fd_sc_hd__a22o_1 _08810_ (.A1(\r1.regblock[0][26] ),
    .A2(_04708_),
    .B1(_04715_),
    .B2(_04712_),
    .X(_03223_));
 sky130_fd_sc_hd__clkbuf_1 _08811_ (.A(_04714_),
    .X(_02197_));
 sky130_fd_sc_hd__buf_1 _08812_ (.A(_04707_),
    .X(_04716_));
 sky130_fd_sc_hd__buf_1 _08813_ (.A(_04485_),
    .X(_04717_));
 sky130_fd_sc_hd__buf_1 _08814_ (.A(_04711_),
    .X(_04718_));
 sky130_fd_sc_hd__a22o_1 _08815_ (.A1(\r1.regblock[0][25] ),
    .A2(_04716_),
    .B1(_04717_),
    .B2(_04718_),
    .X(_03222_));
 sky130_fd_sc_hd__clkbuf_1 _08816_ (.A(_04714_),
    .X(_02196_));
 sky130_fd_sc_hd__buf_1 _08817_ (.A(_04489_),
    .X(_04719_));
 sky130_fd_sc_hd__a22o_1 _08818_ (.A1(\r1.regblock[0][24] ),
    .A2(_04716_),
    .B1(_04719_),
    .B2(_04718_),
    .X(_03221_));
 sky130_fd_sc_hd__buf_2 _08819_ (.A(_04691_),
    .X(_04720_));
 sky130_fd_sc_hd__clkbuf_2 _08820_ (.A(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__clkbuf_1 _08821_ (.A(_04721_),
    .X(_02195_));
 sky130_fd_sc_hd__buf_1 _08822_ (.A(_04493_),
    .X(_04722_));
 sky130_fd_sc_hd__a22o_1 _08823_ (.A1(\r1.regblock[0][23] ),
    .A2(_04716_),
    .B1(_04722_),
    .B2(_04718_),
    .X(_03220_));
 sky130_fd_sc_hd__clkbuf_1 _08824_ (.A(_04721_),
    .X(_02194_));
 sky130_fd_sc_hd__buf_1 _08825_ (.A(_04707_),
    .X(_04723_));
 sky130_fd_sc_hd__buf_1 _08826_ (.A(_04497_),
    .X(_04724_));
 sky130_fd_sc_hd__buf_1 _08827_ (.A(_04711_),
    .X(_04725_));
 sky130_fd_sc_hd__a22o_1 _08828_ (.A1(\r1.regblock[0][22] ),
    .A2(_04723_),
    .B1(_04724_),
    .B2(_04725_),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_1 _08829_ (.A(_04721_),
    .X(_02193_));
 sky130_fd_sc_hd__buf_1 _08830_ (.A(_04501_),
    .X(_04726_));
 sky130_fd_sc_hd__a22o_1 _08831_ (.A1(\r1.regblock[0][21] ),
    .A2(_04723_),
    .B1(_04726_),
    .B2(_04725_),
    .X(_03218_));
 sky130_fd_sc_hd__buf_2 _08832_ (.A(_04720_),
    .X(_04727_));
 sky130_fd_sc_hd__clkbuf_1 _08833_ (.A(_04727_),
    .X(_02192_));
 sky130_fd_sc_hd__buf_1 _08834_ (.A(_04505_),
    .X(_04728_));
 sky130_fd_sc_hd__a22o_1 _08835_ (.A1(\r1.regblock[0][20] ),
    .A2(_04723_),
    .B1(_04728_),
    .B2(_04725_),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_1 _08836_ (.A(_04727_),
    .X(_02191_));
 sky130_fd_sc_hd__clkbuf_2 _08837_ (.A(_04706_),
    .X(_04729_));
 sky130_fd_sc_hd__buf_1 _08838_ (.A(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__buf_1 _08839_ (.A(_04510_),
    .X(_04731_));
 sky130_fd_sc_hd__clkbuf_2 _08840_ (.A(_04710_),
    .X(_04732_));
 sky130_fd_sc_hd__buf_1 _08841_ (.A(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__a22o_1 _08842_ (.A1(\r1.regblock[0][19] ),
    .A2(_04730_),
    .B1(_04731_),
    .B2(_04733_),
    .X(_03216_));
 sky130_fd_sc_hd__clkbuf_1 _08843_ (.A(_04727_),
    .X(_02190_));
 sky130_fd_sc_hd__buf_1 _08844_ (.A(_04515_),
    .X(_04734_));
 sky130_fd_sc_hd__a22o_1 _08845_ (.A1(\r1.regblock[0][18] ),
    .A2(_04730_),
    .B1(_04734_),
    .B2(_04733_),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_2 _08846_ (.A(_04720_),
    .X(_04735_));
 sky130_fd_sc_hd__clkbuf_1 _08847_ (.A(_04735_),
    .X(_02189_));
 sky130_fd_sc_hd__buf_1 _08848_ (.A(_04521_),
    .X(_04736_));
 sky130_fd_sc_hd__a22o_1 _08849_ (.A1(\r1.regblock[0][17] ),
    .A2(_04730_),
    .B1(_04736_),
    .B2(_04733_),
    .X(_03214_));
 sky130_fd_sc_hd__clkbuf_1 _08850_ (.A(_04735_),
    .X(_02188_));
 sky130_fd_sc_hd__buf_1 _08851_ (.A(_04729_),
    .X(_04737_));
 sky130_fd_sc_hd__buf_1 _08852_ (.A(_04525_),
    .X(_04738_));
 sky130_fd_sc_hd__buf_1 _08853_ (.A(_04732_),
    .X(_04739_));
 sky130_fd_sc_hd__a22o_1 _08854_ (.A1(\r1.regblock[0][16] ),
    .A2(_04737_),
    .B1(_04738_),
    .B2(_04739_),
    .X(_03213_));
 sky130_fd_sc_hd__clkbuf_1 _08855_ (.A(_04735_),
    .X(_02187_));
 sky130_fd_sc_hd__buf_1 _08856_ (.A(_04529_),
    .X(_04740_));
 sky130_fd_sc_hd__a22o_1 _08857_ (.A1(\r1.regblock[0][15] ),
    .A2(_04737_),
    .B1(_04740_),
    .B2(_04739_),
    .X(_03212_));
 sky130_fd_sc_hd__buf_2 _08858_ (.A(_04691_),
    .X(_04741_));
 sky130_fd_sc_hd__buf_1 _08859_ (.A(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__clkbuf_1 _08860_ (.A(_04742_),
    .X(_02186_));
 sky130_fd_sc_hd__buf_1 _08861_ (.A(_04533_),
    .X(_04743_));
 sky130_fd_sc_hd__a22o_1 _08862_ (.A1(\r1.regblock[0][14] ),
    .A2(_04737_),
    .B1(_04743_),
    .B2(_04739_),
    .X(_03211_));
 sky130_fd_sc_hd__clkbuf_1 _08863_ (.A(_04742_),
    .X(_02185_));
 sky130_fd_sc_hd__buf_1 _08864_ (.A(_04729_),
    .X(_04744_));
 sky130_fd_sc_hd__buf_1 _08865_ (.A(_04537_),
    .X(_04745_));
 sky130_fd_sc_hd__buf_1 _08866_ (.A(_04732_),
    .X(_04746_));
 sky130_fd_sc_hd__a22o_1 _08867_ (.A1(\r1.regblock[0][13] ),
    .A2(_04744_),
    .B1(_04745_),
    .B2(_04746_),
    .X(_03210_));
 sky130_fd_sc_hd__clkbuf_1 _08868_ (.A(_04742_),
    .X(_02184_));
 sky130_fd_sc_hd__buf_1 _08869_ (.A(_04541_),
    .X(_04747_));
 sky130_fd_sc_hd__a22o_1 _08870_ (.A1(\r1.regblock[0][12] ),
    .A2(_04744_),
    .B1(_04747_),
    .B2(_04746_),
    .X(_03209_));
 sky130_fd_sc_hd__buf_2 _08871_ (.A(_04741_),
    .X(_04748_));
 sky130_fd_sc_hd__clkbuf_1 _08872_ (.A(_04748_),
    .X(_02183_));
 sky130_fd_sc_hd__buf_1 _08873_ (.A(_04545_),
    .X(_04749_));
 sky130_fd_sc_hd__a22o_1 _08874_ (.A1(\r1.regblock[0][11] ),
    .A2(_04744_),
    .B1(_04749_),
    .B2(_04746_),
    .X(_03208_));
 sky130_fd_sc_hd__clkbuf_1 _08875_ (.A(_04748_),
    .X(_02182_));
 sky130_fd_sc_hd__buf_1 _08876_ (.A(_04706_),
    .X(_04750_));
 sky130_fd_sc_hd__buf_1 _08877_ (.A(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__buf_1 _08878_ (.A(_04550_),
    .X(_04752_));
 sky130_fd_sc_hd__buf_1 _08879_ (.A(_04710_),
    .X(_04753_));
 sky130_fd_sc_hd__buf_1 _08880_ (.A(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__a22o_1 _08881_ (.A1(\r1.regblock[0][10] ),
    .A2(_04751_),
    .B1(_04752_),
    .B2(_04754_),
    .X(_03207_));
 sky130_fd_sc_hd__clkbuf_1 _08882_ (.A(_04748_),
    .X(_02181_));
 sky130_fd_sc_hd__buf_1 _08883_ (.A(_04555_),
    .X(_04755_));
 sky130_fd_sc_hd__a22o_1 _08884_ (.A1(\r1.regblock[0][9] ),
    .A2(_04751_),
    .B1(_04755_),
    .B2(_04754_),
    .X(_03206_));
 sky130_fd_sc_hd__buf_1 _08885_ (.A(_04741_),
    .X(_04756_));
 sky130_fd_sc_hd__clkbuf_1 _08886_ (.A(_04756_),
    .X(_02180_));
 sky130_fd_sc_hd__buf_1 _08887_ (.A(_04560_),
    .X(_04757_));
 sky130_fd_sc_hd__a22o_1 _08888_ (.A1(\r1.regblock[0][8] ),
    .A2(_04751_),
    .B1(_04757_),
    .B2(_04754_),
    .X(_03205_));
 sky130_fd_sc_hd__clkbuf_1 _08889_ (.A(_04756_),
    .X(_02179_));
 sky130_fd_sc_hd__buf_1 _08890_ (.A(_04750_),
    .X(_04758_));
 sky130_fd_sc_hd__buf_1 _08891_ (.A(_04564_),
    .X(_04759_));
 sky130_fd_sc_hd__buf_1 _08892_ (.A(_04753_),
    .X(_04760_));
 sky130_fd_sc_hd__a22o_1 _08893_ (.A1(\r1.regblock[0][7] ),
    .A2(_04758_),
    .B1(_04759_),
    .B2(_04760_),
    .X(_03204_));
 sky130_fd_sc_hd__clkbuf_1 _08894_ (.A(_04756_),
    .X(_02178_));
 sky130_fd_sc_hd__buf_1 _08895_ (.A(_04568_),
    .X(_04761_));
 sky130_fd_sc_hd__a22o_1 _08896_ (.A1(\r1.regblock[0][6] ),
    .A2(_04758_),
    .B1(_04761_),
    .B2(_04760_),
    .X(_03203_));
 sky130_fd_sc_hd__buf_2 _08897_ (.A(_04657_),
    .X(_04762_));
 sky130_fd_sc_hd__clkbuf_2 _08898_ (.A(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__buf_1 _08899_ (.A(_04763_),
    .X(_04764_));
 sky130_fd_sc_hd__clkbuf_1 _08900_ (.A(_04764_),
    .X(_02177_));
 sky130_fd_sc_hd__buf_1 _08901_ (.A(_04572_),
    .X(_04765_));
 sky130_fd_sc_hd__a22o_1 _08902_ (.A1(\r1.regblock[0][5] ),
    .A2(_04758_),
    .B1(_04765_),
    .B2(_04760_),
    .X(_03202_));
 sky130_fd_sc_hd__clkbuf_1 _08903_ (.A(_04764_),
    .X(_02176_));
 sky130_fd_sc_hd__buf_1 _08904_ (.A(_04750_),
    .X(_04766_));
 sky130_fd_sc_hd__buf_1 _08905_ (.A(_04576_),
    .X(_04767_));
 sky130_fd_sc_hd__buf_1 _08906_ (.A(_04753_),
    .X(_04768_));
 sky130_fd_sc_hd__a22o_1 _08907_ (.A1(\r1.regblock[0][4] ),
    .A2(_04766_),
    .B1(_04767_),
    .B2(_04768_),
    .X(_03201_));
 sky130_fd_sc_hd__clkbuf_1 _08908_ (.A(_04764_),
    .X(_02175_));
 sky130_fd_sc_hd__buf_1 _08909_ (.A(_04580_),
    .X(_04769_));
 sky130_fd_sc_hd__a22o_1 _08910_ (.A1(\r1.regblock[0][3] ),
    .A2(_04766_),
    .B1(_04769_),
    .B2(_04768_),
    .X(_03200_));
 sky130_fd_sc_hd__clkbuf_2 _08911_ (.A(_04763_),
    .X(_04770_));
 sky130_fd_sc_hd__clkbuf_1 _08912_ (.A(_04770_),
    .X(_02174_));
 sky130_fd_sc_hd__buf_1 _08913_ (.A(_04584_),
    .X(_04771_));
 sky130_fd_sc_hd__a22o_1 _08914_ (.A1(\r1.regblock[0][2] ),
    .A2(_04766_),
    .B1(_04771_),
    .B2(_04768_),
    .X(_03199_));
 sky130_fd_sc_hd__clkbuf_1 _08915_ (.A(_04770_),
    .X(_02173_));
 sky130_fd_sc_hd__buf_1 _08916_ (.A(_04587_),
    .X(_04772_));
 sky130_fd_sc_hd__a22o_1 _08917_ (.A1(\r1.regblock[0][1] ),
    .A2(_04697_),
    .B1(_04772_),
    .B2(_04701_),
    .X(_03198_));
 sky130_fd_sc_hd__clkbuf_1 _08918_ (.A(_04770_),
    .X(_02172_));
 sky130_fd_sc_hd__buf_1 _08919_ (.A(_04590_),
    .X(_04773_));
 sky130_fd_sc_hd__a22o_1 _08920_ (.A1(\r1.regblock[0][0] ),
    .A2(_04697_),
    .B1(_04773_),
    .B2(_04701_),
    .X(_03197_));
 sky130_fd_sc_hd__buf_1 _08921_ (.A(_04763_),
    .X(_04774_));
 sky130_fd_sc_hd__clkbuf_1 _08922_ (.A(_04774_),
    .X(_02171_));
 sky130_fd_sc_hd__buf_1 _08923_ (.A(_04694_),
    .X(_04775_));
 sky130_fd_sc_hd__buf_1 _08924_ (.A(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__or3_1 _08925_ (.A(_04213_),
    .B(_04390_),
    .C(_04215_),
    .X(_04777_));
 sky130_fd_sc_hd__clkbuf_1 _08926_ (.A(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__or2_2 _08927_ (.A(_04776_),
    .B(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__buf_1 _08928_ (.A(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__buf_1 _08929_ (.A(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__inv_2 _08930_ (.A(_04779_),
    .Y(_04782_));
 sky130_fd_sc_hd__buf_1 _08931_ (.A(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__buf_1 _08932_ (.A(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__a22o_1 _08933_ (.A1(\r1.regblock[8][31] ),
    .A2(_04781_),
    .B1(_04699_),
    .B2(_04784_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_1 _08934_ (.A(_04774_),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_1 _08935_ (.A1(\r1.regblock[8][30] ),
    .A2(_04781_),
    .B1(_04703_),
    .B2(_04784_),
    .X(_03195_));
 sky130_fd_sc_hd__clkbuf_1 _08936_ (.A(_04774_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _08937_ (.A1(\r1.regblock[8][29] ),
    .A2(_04781_),
    .B1(_04705_),
    .B2(_04784_),
    .X(_03194_));
 sky130_fd_sc_hd__clkbuf_2 _08938_ (.A(_04762_),
    .X(_04785_));
 sky130_fd_sc_hd__buf_1 _08939_ (.A(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__clkbuf_1 _08940_ (.A(_04786_),
    .X(_02168_));
 sky130_fd_sc_hd__clkbuf_4 _08941_ (.A(_04779_),
    .X(_04787_));
 sky130_fd_sc_hd__clkbuf_2 _08942_ (.A(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__buf_1 _08943_ (.A(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__clkbuf_4 _08944_ (.A(_04782_),
    .X(_04790_));
 sky130_fd_sc_hd__clkbuf_2 _08945_ (.A(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__buf_1 _08946_ (.A(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__a22o_1 _08947_ (.A1(\r1.regblock[8][28] ),
    .A2(_04789_),
    .B1(_04709_),
    .B2(_04792_),
    .X(_03193_));
 sky130_fd_sc_hd__clkbuf_1 _08948_ (.A(_04786_),
    .X(_02167_));
 sky130_fd_sc_hd__a22o_1 _08949_ (.A1(\r1.regblock[8][27] ),
    .A2(_04789_),
    .B1(_04713_),
    .B2(_04792_),
    .X(_03192_));
 sky130_fd_sc_hd__clkbuf_1 _08950_ (.A(_04786_),
    .X(_02166_));
 sky130_fd_sc_hd__a22o_1 _08951_ (.A1(\r1.regblock[8][26] ),
    .A2(_04789_),
    .B1(_04715_),
    .B2(_04792_),
    .X(_03191_));
 sky130_fd_sc_hd__buf_1 _08952_ (.A(_04785_),
    .X(_04793_));
 sky130_fd_sc_hd__clkbuf_1 _08953_ (.A(_04793_),
    .X(_02165_));
 sky130_fd_sc_hd__buf_1 _08954_ (.A(_04788_),
    .X(_04794_));
 sky130_fd_sc_hd__buf_1 _08955_ (.A(_04791_),
    .X(_04795_));
 sky130_fd_sc_hd__a22o_1 _08956_ (.A1(\r1.regblock[8][25] ),
    .A2(_04794_),
    .B1(_04717_),
    .B2(_04795_),
    .X(_03190_));
 sky130_fd_sc_hd__clkbuf_1 _08957_ (.A(_04793_),
    .X(_02164_));
 sky130_fd_sc_hd__a22o_1 _08958_ (.A1(\r1.regblock[8][24] ),
    .A2(_04794_),
    .B1(_04719_),
    .B2(_04795_),
    .X(_03189_));
 sky130_fd_sc_hd__clkbuf_1 _08959_ (.A(_04793_),
    .X(_02163_));
 sky130_fd_sc_hd__a22o_1 _08960_ (.A1(\r1.regblock[8][23] ),
    .A2(_04794_),
    .B1(_04722_),
    .B2(_04795_),
    .X(_03188_));
 sky130_fd_sc_hd__buf_1 _08961_ (.A(_04785_),
    .X(_04796_));
 sky130_fd_sc_hd__clkbuf_1 _08962_ (.A(_04796_),
    .X(_02162_));
 sky130_fd_sc_hd__buf_1 _08963_ (.A(_04788_),
    .X(_04797_));
 sky130_fd_sc_hd__buf_1 _08964_ (.A(_04791_),
    .X(_04798_));
 sky130_fd_sc_hd__a22o_1 _08965_ (.A1(\r1.regblock[8][22] ),
    .A2(_04797_),
    .B1(_04724_),
    .B2(_04798_),
    .X(_03187_));
 sky130_fd_sc_hd__clkbuf_1 _08966_ (.A(_04796_),
    .X(_02161_));
 sky130_fd_sc_hd__a22o_1 _08967_ (.A1(\r1.regblock[8][21] ),
    .A2(_04797_),
    .B1(_04726_),
    .B2(_04798_),
    .X(_03186_));
 sky130_fd_sc_hd__clkbuf_1 _08968_ (.A(_04796_),
    .X(_02160_));
 sky130_fd_sc_hd__a22o_1 _08969_ (.A1(\r1.regblock[8][20] ),
    .A2(_04797_),
    .B1(_04728_),
    .B2(_04798_),
    .X(_03185_));
 sky130_fd_sc_hd__clkbuf_2 _08970_ (.A(_04762_),
    .X(_04799_));
 sky130_fd_sc_hd__buf_1 _08971_ (.A(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__clkbuf_1 _08972_ (.A(_04800_),
    .X(_02159_));
 sky130_fd_sc_hd__clkbuf_2 _08973_ (.A(_04787_),
    .X(_04801_));
 sky130_fd_sc_hd__buf_1 _08974_ (.A(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__buf_2 _08975_ (.A(_04790_),
    .X(_04803_));
 sky130_fd_sc_hd__buf_1 _08976_ (.A(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__a22o_1 _08977_ (.A1(\r1.regblock[8][19] ),
    .A2(_04802_),
    .B1(_04731_),
    .B2(_04804_),
    .X(_03184_));
 sky130_fd_sc_hd__clkbuf_1 _08978_ (.A(_04800_),
    .X(_02158_));
 sky130_fd_sc_hd__a22o_1 _08979_ (.A1(\r1.regblock[8][18] ),
    .A2(_04802_),
    .B1(_04734_),
    .B2(_04804_),
    .X(_03183_));
 sky130_fd_sc_hd__clkbuf_1 _08980_ (.A(_04800_),
    .X(_02157_));
 sky130_fd_sc_hd__a22o_1 _08981_ (.A1(\r1.regblock[8][17] ),
    .A2(_04802_),
    .B1(_04736_),
    .B2(_04804_),
    .X(_03182_));
 sky130_fd_sc_hd__buf_1 _08982_ (.A(_04799_),
    .X(_04805_));
 sky130_fd_sc_hd__clkbuf_1 _08983_ (.A(_04805_),
    .X(_02156_));
 sky130_fd_sc_hd__buf_1 _08984_ (.A(_04801_),
    .X(_04806_));
 sky130_fd_sc_hd__buf_1 _08985_ (.A(_04803_),
    .X(_04807_));
 sky130_fd_sc_hd__a22o_1 _08986_ (.A1(\r1.regblock[8][16] ),
    .A2(_04806_),
    .B1(_04738_),
    .B2(_04807_),
    .X(_03181_));
 sky130_fd_sc_hd__clkbuf_1 _08987_ (.A(_04805_),
    .X(_02155_));
 sky130_fd_sc_hd__a22o_1 _08988_ (.A1(\r1.regblock[8][15] ),
    .A2(_04806_),
    .B1(_04740_),
    .B2(_04807_),
    .X(_03180_));
 sky130_fd_sc_hd__clkbuf_1 _08989_ (.A(_04805_),
    .X(_02154_));
 sky130_fd_sc_hd__a22o_1 _08990_ (.A1(\r1.regblock[8][14] ),
    .A2(_04806_),
    .B1(_04743_),
    .B2(_04807_),
    .X(_03179_));
 sky130_fd_sc_hd__buf_1 _08991_ (.A(_04799_),
    .X(_04808_));
 sky130_fd_sc_hd__clkbuf_1 _08992_ (.A(_04808_),
    .X(_02153_));
 sky130_fd_sc_hd__buf_1 _08993_ (.A(_04801_),
    .X(_04809_));
 sky130_fd_sc_hd__buf_1 _08994_ (.A(_04803_),
    .X(_04810_));
 sky130_fd_sc_hd__a22o_1 _08995_ (.A1(\r1.regblock[8][13] ),
    .A2(_04809_),
    .B1(_04745_),
    .B2(_04810_),
    .X(_03178_));
 sky130_fd_sc_hd__clkbuf_1 _08996_ (.A(_04808_),
    .X(_02152_));
 sky130_fd_sc_hd__a22o_1 _08997_ (.A1(\r1.regblock[8][12] ),
    .A2(_04809_),
    .B1(_04747_),
    .B2(_04810_),
    .X(_03177_));
 sky130_fd_sc_hd__clkbuf_1 _08998_ (.A(_04808_),
    .X(_02151_));
 sky130_fd_sc_hd__a22o_1 _08999_ (.A1(\r1.regblock[8][11] ),
    .A2(_04809_),
    .B1(_04749_),
    .B2(_04810_),
    .X(_03176_));
 sky130_fd_sc_hd__buf_1 _09000_ (.A(_04430_),
    .X(_04811_));
 sky130_fd_sc_hd__buf_1 _09001_ (.A(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__clkbuf_2 _09002_ (.A(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__buf_1 _09003_ (.A(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__clkbuf_1 _09004_ (.A(_04814_),
    .X(_02150_));
 sky130_fd_sc_hd__clkbuf_2 _09005_ (.A(_04787_),
    .X(_04815_));
 sky130_fd_sc_hd__buf_1 _09006_ (.A(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__clkbuf_2 _09007_ (.A(_04790_),
    .X(_04817_));
 sky130_fd_sc_hd__buf_1 _09008_ (.A(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__a22o_1 _09009_ (.A1(\r1.regblock[8][10] ),
    .A2(_04816_),
    .B1(_04752_),
    .B2(_04818_),
    .X(_03175_));
 sky130_fd_sc_hd__clkbuf_1 _09010_ (.A(_04814_),
    .X(_02149_));
 sky130_fd_sc_hd__a22o_1 _09011_ (.A1(\r1.regblock[8][9] ),
    .A2(_04816_),
    .B1(_04755_),
    .B2(_04818_),
    .X(_03174_));
 sky130_fd_sc_hd__clkbuf_1 _09012_ (.A(_04814_),
    .X(_02148_));
 sky130_fd_sc_hd__a22o_1 _09013_ (.A1(\r1.regblock[8][8] ),
    .A2(_04816_),
    .B1(_04757_),
    .B2(_04818_),
    .X(_03173_));
 sky130_fd_sc_hd__buf_1 _09014_ (.A(_04813_),
    .X(_04819_));
 sky130_fd_sc_hd__clkbuf_1 _09015_ (.A(_04819_),
    .X(_02147_));
 sky130_fd_sc_hd__buf_1 _09016_ (.A(_04815_),
    .X(_04820_));
 sky130_fd_sc_hd__buf_1 _09017_ (.A(_04817_),
    .X(_04821_));
 sky130_fd_sc_hd__a22o_1 _09018_ (.A1(\r1.regblock[8][7] ),
    .A2(_04820_),
    .B1(_04759_),
    .B2(_04821_),
    .X(_03172_));
 sky130_fd_sc_hd__clkbuf_1 _09019_ (.A(_04819_),
    .X(_02146_));
 sky130_fd_sc_hd__a22o_1 _09020_ (.A1(\r1.regblock[8][6] ),
    .A2(_04820_),
    .B1(_04761_),
    .B2(_04821_),
    .X(_03171_));
 sky130_fd_sc_hd__clkbuf_1 _09021_ (.A(_04819_),
    .X(_02145_));
 sky130_fd_sc_hd__a22o_1 _09022_ (.A1(\r1.regblock[8][5] ),
    .A2(_04820_),
    .B1(_04765_),
    .B2(_04821_),
    .X(_03170_));
 sky130_fd_sc_hd__buf_1 _09023_ (.A(_04813_),
    .X(_04822_));
 sky130_fd_sc_hd__clkbuf_1 _09024_ (.A(_04822_),
    .X(_02144_));
 sky130_fd_sc_hd__buf_1 _09025_ (.A(_04815_),
    .X(_04823_));
 sky130_fd_sc_hd__buf_1 _09026_ (.A(_04817_),
    .X(_04824_));
 sky130_fd_sc_hd__a22o_1 _09027_ (.A1(\r1.regblock[8][4] ),
    .A2(_04823_),
    .B1(_04767_),
    .B2(_04824_),
    .X(_03169_));
 sky130_fd_sc_hd__clkbuf_1 _09028_ (.A(_04822_),
    .X(_02143_));
 sky130_fd_sc_hd__a22o_1 _09029_ (.A1(\r1.regblock[8][3] ),
    .A2(_04823_),
    .B1(_04769_),
    .B2(_04824_),
    .X(_03168_));
 sky130_fd_sc_hd__clkbuf_1 _09030_ (.A(_04822_),
    .X(_02142_));
 sky130_fd_sc_hd__a22o_1 _09031_ (.A1(\r1.regblock[8][2] ),
    .A2(_04823_),
    .B1(_04771_),
    .B2(_04824_),
    .X(_03167_));
 sky130_fd_sc_hd__buf_2 _09032_ (.A(_04812_),
    .X(_04825_));
 sky130_fd_sc_hd__buf_1 _09033_ (.A(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__clkbuf_1 _09034_ (.A(_04826_),
    .X(_02141_));
 sky130_fd_sc_hd__a22o_1 _09035_ (.A1(\r1.regblock[8][1] ),
    .A2(_04780_),
    .B1(_04772_),
    .B2(_04783_),
    .X(_03166_));
 sky130_fd_sc_hd__clkbuf_1 _09036_ (.A(_04826_),
    .X(_02140_));
 sky130_fd_sc_hd__a22o_1 _09037_ (.A1(\r1.regblock[8][0] ),
    .A2(_04780_),
    .B1(_04773_),
    .B2(_04783_),
    .X(_03165_));
 sky130_fd_sc_hd__clkbuf_1 _09038_ (.A(_04826_),
    .X(_02139_));
 sky130_fd_sc_hd__or2_2 _09039_ (.A(_04641_),
    .B(_04778_),
    .X(_04827_));
 sky130_fd_sc_hd__buf_1 _09040_ (.A(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__buf_1 _09041_ (.A(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__inv_2 _09042_ (.A(_04827_),
    .Y(_04830_));
 sky130_fd_sc_hd__buf_1 _09043_ (.A(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__buf_1 _09044_ (.A(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__a22o_1 _09045_ (.A1(\r1.regblock[9][31] ),
    .A2(_04829_),
    .B1(_04699_),
    .B2(_04832_),
    .X(_03164_));
 sky130_fd_sc_hd__clkbuf_2 _09046_ (.A(_04825_),
    .X(_04833_));
 sky130_fd_sc_hd__clkbuf_1 _09047_ (.A(_04833_),
    .X(_02138_));
 sky130_fd_sc_hd__a22o_1 _09048_ (.A1(\r1.regblock[9][30] ),
    .A2(_04829_),
    .B1(_04703_),
    .B2(_04832_),
    .X(_03163_));
 sky130_fd_sc_hd__clkbuf_1 _09049_ (.A(_04833_),
    .X(_02137_));
 sky130_fd_sc_hd__a22o_1 _09050_ (.A1(\r1.regblock[9][29] ),
    .A2(_04829_),
    .B1(_04705_),
    .B2(_04832_),
    .X(_03162_));
 sky130_fd_sc_hd__clkbuf_1 _09051_ (.A(_04833_),
    .X(_02136_));
 sky130_fd_sc_hd__clkbuf_4 _09052_ (.A(_04827_),
    .X(_04834_));
 sky130_fd_sc_hd__clkbuf_2 _09053_ (.A(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__buf_1 _09054_ (.A(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__clkbuf_4 _09055_ (.A(_04830_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_2 _09056_ (.A(_04837_),
    .X(_04838_));
 sky130_fd_sc_hd__buf_1 _09057_ (.A(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__a22o_1 _09058_ (.A1(\r1.regblock[9][28] ),
    .A2(_04836_),
    .B1(_04709_),
    .B2(_04839_),
    .X(_03161_));
 sky130_fd_sc_hd__buf_1 _09059_ (.A(_04825_),
    .X(_04840_));
 sky130_fd_sc_hd__clkbuf_1 _09060_ (.A(_04840_),
    .X(_02135_));
 sky130_fd_sc_hd__a22o_1 _09061_ (.A1(\r1.regblock[9][27] ),
    .A2(_04836_),
    .B1(_04713_),
    .B2(_04839_),
    .X(_03160_));
 sky130_fd_sc_hd__clkbuf_1 _09062_ (.A(_04840_),
    .X(_02134_));
 sky130_fd_sc_hd__a22o_1 _09063_ (.A1(\r1.regblock[9][26] ),
    .A2(_04836_),
    .B1(_04715_),
    .B2(_04839_),
    .X(_03159_));
 sky130_fd_sc_hd__clkbuf_1 _09064_ (.A(_04840_),
    .X(_02133_));
 sky130_fd_sc_hd__buf_1 _09065_ (.A(_04835_),
    .X(_04841_));
 sky130_fd_sc_hd__buf_1 _09066_ (.A(_04838_),
    .X(_04842_));
 sky130_fd_sc_hd__a22o_1 _09067_ (.A1(\r1.regblock[9][25] ),
    .A2(_04841_),
    .B1(_04717_),
    .B2(_04842_),
    .X(_03158_));
 sky130_fd_sc_hd__buf_2 _09068_ (.A(_04812_),
    .X(_04843_));
 sky130_fd_sc_hd__buf_1 _09069_ (.A(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__clkbuf_1 _09070_ (.A(_04844_),
    .X(_02132_));
 sky130_fd_sc_hd__a22o_1 _09071_ (.A1(\r1.regblock[9][24] ),
    .A2(_04841_),
    .B1(_04719_),
    .B2(_04842_),
    .X(_03157_));
 sky130_fd_sc_hd__clkbuf_1 _09072_ (.A(_04844_),
    .X(_02131_));
 sky130_fd_sc_hd__a22o_1 _09073_ (.A1(\r1.regblock[9][23] ),
    .A2(_04841_),
    .B1(_04722_),
    .B2(_04842_),
    .X(_03156_));
 sky130_fd_sc_hd__clkbuf_1 _09074_ (.A(_04844_),
    .X(_02130_));
 sky130_fd_sc_hd__buf_1 _09075_ (.A(_04835_),
    .X(_04845_));
 sky130_fd_sc_hd__buf_1 _09076_ (.A(_04838_),
    .X(_04846_));
 sky130_fd_sc_hd__a22o_1 _09077_ (.A1(\r1.regblock[9][22] ),
    .A2(_04845_),
    .B1(_04724_),
    .B2(_04846_),
    .X(_03155_));
 sky130_fd_sc_hd__buf_2 _09078_ (.A(_04843_),
    .X(_04847_));
 sky130_fd_sc_hd__clkbuf_1 _09079_ (.A(_04847_),
    .X(_02129_));
 sky130_fd_sc_hd__a22o_1 _09080_ (.A1(\r1.regblock[9][21] ),
    .A2(_04845_),
    .B1(_04726_),
    .B2(_04846_),
    .X(_03154_));
 sky130_fd_sc_hd__clkbuf_1 _09081_ (.A(_04847_),
    .X(_02128_));
 sky130_fd_sc_hd__a22o_1 _09082_ (.A1(\r1.regblock[9][20] ),
    .A2(_04845_),
    .B1(_04728_),
    .B2(_04846_),
    .X(_03153_));
 sky130_fd_sc_hd__clkbuf_1 _09083_ (.A(_04847_),
    .X(_02127_));
 sky130_fd_sc_hd__clkbuf_2 _09084_ (.A(_04834_),
    .X(_04848_));
 sky130_fd_sc_hd__buf_1 _09085_ (.A(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__clkbuf_2 _09086_ (.A(_04837_),
    .X(_04850_));
 sky130_fd_sc_hd__buf_1 _09087_ (.A(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__a22o_1 _09088_ (.A1(\r1.regblock[9][19] ),
    .A2(_04849_),
    .B1(_04731_),
    .B2(_04851_),
    .X(_03152_));
 sky130_fd_sc_hd__buf_1 _09089_ (.A(_04843_),
    .X(_04852_));
 sky130_fd_sc_hd__clkbuf_1 _09090_ (.A(_04852_),
    .X(_02126_));
 sky130_fd_sc_hd__a22o_1 _09091_ (.A1(\r1.regblock[9][18] ),
    .A2(_04849_),
    .B1(_04734_),
    .B2(_04851_),
    .X(_03151_));
 sky130_fd_sc_hd__clkbuf_1 _09092_ (.A(_04852_),
    .X(_02125_));
 sky130_fd_sc_hd__a22o_1 _09093_ (.A1(\r1.regblock[9][17] ),
    .A2(_04849_),
    .B1(_04736_),
    .B2(_04851_),
    .X(_03150_));
 sky130_fd_sc_hd__clkbuf_1 _09094_ (.A(_04852_),
    .X(_02124_));
 sky130_fd_sc_hd__buf_1 _09095_ (.A(_04848_),
    .X(_04853_));
 sky130_fd_sc_hd__buf_1 _09096_ (.A(_04850_),
    .X(_04854_));
 sky130_fd_sc_hd__a22o_1 _09097_ (.A1(\r1.regblock[9][16] ),
    .A2(_04853_),
    .B1(_04738_),
    .B2(_04854_),
    .X(_03149_));
 sky130_fd_sc_hd__clkbuf_2 _09098_ (.A(_04811_),
    .X(_04855_));
 sky130_fd_sc_hd__buf_2 _09099_ (.A(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__buf_1 _09100_ (.A(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_1 _09101_ (.A(_04857_),
    .X(_02123_));
 sky130_fd_sc_hd__a22o_1 _09102_ (.A1(\r1.regblock[9][15] ),
    .A2(_04853_),
    .B1(_04740_),
    .B2(_04854_),
    .X(_03148_));
 sky130_fd_sc_hd__clkbuf_1 _09103_ (.A(_04857_),
    .X(_02122_));
 sky130_fd_sc_hd__a22o_1 _09104_ (.A1(\r1.regblock[9][14] ),
    .A2(_04853_),
    .B1(_04743_),
    .B2(_04854_),
    .X(_03147_));
 sky130_fd_sc_hd__clkbuf_1 _09105_ (.A(_04857_),
    .X(_02121_));
 sky130_fd_sc_hd__buf_1 _09106_ (.A(_04848_),
    .X(_04858_));
 sky130_fd_sc_hd__buf_1 _09107_ (.A(_04850_),
    .X(_04859_));
 sky130_fd_sc_hd__a22o_1 _09108_ (.A1(\r1.regblock[9][13] ),
    .A2(_04858_),
    .B1(_04745_),
    .B2(_04859_),
    .X(_03146_));
 sky130_fd_sc_hd__buf_1 _09109_ (.A(_04856_),
    .X(_04860_));
 sky130_fd_sc_hd__clkbuf_1 _09110_ (.A(_04860_),
    .X(_02120_));
 sky130_fd_sc_hd__a22o_1 _09111_ (.A1(\r1.regblock[9][12] ),
    .A2(_04858_),
    .B1(_04747_),
    .B2(_04859_),
    .X(_03145_));
 sky130_fd_sc_hd__clkbuf_1 _09112_ (.A(_04860_),
    .X(_02119_));
 sky130_fd_sc_hd__a22o_1 _09113_ (.A1(\r1.regblock[9][11] ),
    .A2(_04858_),
    .B1(_04749_),
    .B2(_04859_),
    .X(_03144_));
 sky130_fd_sc_hd__clkbuf_2 _09114_ (.A(_04860_),
    .X(_02118_));
 sky130_fd_sc_hd__buf_1 _09115_ (.A(_04834_),
    .X(_04861_));
 sky130_fd_sc_hd__buf_1 _09116_ (.A(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__buf_1 _09117_ (.A(_04837_),
    .X(_04863_));
 sky130_fd_sc_hd__buf_1 _09118_ (.A(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__a22o_1 _09119_ (.A1(\r1.regblock[9][10] ),
    .A2(_04862_),
    .B1(_04752_),
    .B2(_04864_),
    .X(_03143_));
 sky130_fd_sc_hd__buf_1 _09120_ (.A(_04856_),
    .X(_04865_));
 sky130_fd_sc_hd__clkbuf_1 _09121_ (.A(_04865_),
    .X(_02117_));
 sky130_fd_sc_hd__a22o_1 _09122_ (.A1(\r1.regblock[9][9] ),
    .A2(_04862_),
    .B1(_04755_),
    .B2(_04864_),
    .X(_03142_));
 sky130_fd_sc_hd__clkbuf_1 _09123_ (.A(_04865_),
    .X(_02116_));
 sky130_fd_sc_hd__a22o_1 _09124_ (.A1(\r1.regblock[9][8] ),
    .A2(_04862_),
    .B1(_04757_),
    .B2(_04864_),
    .X(_03141_));
 sky130_fd_sc_hd__clkbuf_1 _09125_ (.A(_04865_),
    .X(_02115_));
 sky130_fd_sc_hd__buf_1 _09126_ (.A(_04861_),
    .X(_04866_));
 sky130_fd_sc_hd__buf_1 _09127_ (.A(_04863_),
    .X(_04867_));
 sky130_fd_sc_hd__a22o_1 _09128_ (.A1(\r1.regblock[9][7] ),
    .A2(_04866_),
    .B1(_04759_),
    .B2(_04867_),
    .X(_03140_));
 sky130_fd_sc_hd__buf_1 _09129_ (.A(_04855_),
    .X(_04868_));
 sky130_fd_sc_hd__buf_1 _09130_ (.A(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__clkbuf_1 _09131_ (.A(_04869_),
    .X(_02114_));
 sky130_fd_sc_hd__a22o_1 _09132_ (.A1(\r1.regblock[9][6] ),
    .A2(_04866_),
    .B1(_04761_),
    .B2(_04867_),
    .X(_03139_));
 sky130_fd_sc_hd__clkbuf_1 _09133_ (.A(_04869_),
    .X(_02113_));
 sky130_fd_sc_hd__a22o_1 _09134_ (.A1(\r1.regblock[9][5] ),
    .A2(_04866_),
    .B1(_04765_),
    .B2(_04867_),
    .X(_03138_));
 sky130_fd_sc_hd__clkbuf_1 _09135_ (.A(_04869_),
    .X(_02112_));
 sky130_fd_sc_hd__buf_1 _09136_ (.A(_04861_),
    .X(_04870_));
 sky130_fd_sc_hd__buf_1 _09137_ (.A(_04863_),
    .X(_04871_));
 sky130_fd_sc_hd__a22o_1 _09138_ (.A1(\r1.regblock[9][4] ),
    .A2(_04870_),
    .B1(_04767_),
    .B2(_04871_),
    .X(_03137_));
 sky130_fd_sc_hd__clkbuf_2 _09139_ (.A(_04868_),
    .X(_04872_));
 sky130_fd_sc_hd__clkbuf_1 _09140_ (.A(_04872_),
    .X(_02111_));
 sky130_fd_sc_hd__a22o_1 _09141_ (.A1(\r1.regblock[9][3] ),
    .A2(_04870_),
    .B1(_04769_),
    .B2(_04871_),
    .X(_03136_));
 sky130_fd_sc_hd__clkbuf_1 _09142_ (.A(_04872_),
    .X(_02110_));
 sky130_fd_sc_hd__a22o_1 _09143_ (.A1(\r1.regblock[9][2] ),
    .A2(_04870_),
    .B1(_04771_),
    .B2(_04871_),
    .X(_03135_));
 sky130_fd_sc_hd__clkbuf_1 _09144_ (.A(_04872_),
    .X(_02109_));
 sky130_fd_sc_hd__a22o_1 _09145_ (.A1(\r1.regblock[9][1] ),
    .A2(_04828_),
    .B1(_04772_),
    .B2(_04831_),
    .X(_03134_));
 sky130_fd_sc_hd__clkbuf_2 _09146_ (.A(_04868_),
    .X(_04873_));
 sky130_fd_sc_hd__clkbuf_1 _09147_ (.A(_04873_),
    .X(_02108_));
 sky130_fd_sc_hd__a22o_1 _09148_ (.A1(\r1.regblock[9][0] ),
    .A2(_04828_),
    .B1(_04773_),
    .B2(_04831_),
    .X(_03133_));
 sky130_fd_sc_hd__clkbuf_1 _09149_ (.A(_04873_),
    .X(_02107_));
 sky130_fd_sc_hd__or2_1 _09150_ (.A(_04394_),
    .B(_04695_),
    .X(_04874_));
 sky130_fd_sc_hd__buf_1 _09151_ (.A(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__buf_1 _09152_ (.A(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__buf_1 _09153_ (.A(_04454_),
    .X(_04877_));
 sky130_fd_sc_hd__inv_2 _09154_ (.A(_04874_),
    .Y(_04878_));
 sky130_fd_sc_hd__buf_1 _09155_ (.A(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__buf_1 _09156_ (.A(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__a22o_1 _09157_ (.A1(\r1.regblock[12][31] ),
    .A2(_04876_),
    .B1(_04877_),
    .B2(_04880_),
    .X(_03132_));
 sky130_fd_sc_hd__clkbuf_1 _09158_ (.A(_04873_),
    .X(_02106_));
 sky130_fd_sc_hd__buf_1 _09159_ (.A(_04460_),
    .X(_04881_));
 sky130_fd_sc_hd__a22o_1 _09160_ (.A1(\r1.regblock[12][30] ),
    .A2(_04876_),
    .B1(_04881_),
    .B2(_04880_),
    .X(_03131_));
 sky130_fd_sc_hd__clkbuf_2 _09161_ (.A(_04855_),
    .X(_04882_));
 sky130_fd_sc_hd__buf_1 _09162_ (.A(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__buf_1 _09163_ (.A(_04883_),
    .X(_02105_));
 sky130_fd_sc_hd__buf_1 _09164_ (.A(_04464_),
    .X(_04884_));
 sky130_fd_sc_hd__a22o_1 _09165_ (.A1(\r1.regblock[12][29] ),
    .A2(_04876_),
    .B1(_04884_),
    .B2(_04880_),
    .X(_03130_));
 sky130_fd_sc_hd__clkbuf_1 _09166_ (.A(_04883_),
    .X(_02104_));
 sky130_fd_sc_hd__buf_2 _09167_ (.A(_04874_),
    .X(_04885_));
 sky130_fd_sc_hd__buf_2 _09168_ (.A(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__buf_1 _09169_ (.A(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__buf_1 _09170_ (.A(_04470_),
    .X(_04888_));
 sky130_fd_sc_hd__buf_2 _09171_ (.A(_04878_),
    .X(_04889_));
 sky130_fd_sc_hd__buf_2 _09172_ (.A(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__buf_1 _09173_ (.A(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__a22o_1 _09174_ (.A1(\r1.regblock[12][28] ),
    .A2(_04887_),
    .B1(_04888_),
    .B2(_04891_),
    .X(_03129_));
 sky130_fd_sc_hd__clkbuf_1 _09175_ (.A(_04883_),
    .X(_02103_));
 sky130_fd_sc_hd__buf_1 _09176_ (.A(_04476_),
    .X(_04892_));
 sky130_fd_sc_hd__a22o_1 _09177_ (.A1(\r1.regblock[12][27] ),
    .A2(_04887_),
    .B1(_04892_),
    .B2(_04891_),
    .X(_03128_));
 sky130_fd_sc_hd__buf_1 _09178_ (.A(_04882_),
    .X(_04893_));
 sky130_fd_sc_hd__buf_1 _09179_ (.A(_04893_),
    .X(_02102_));
 sky130_fd_sc_hd__buf_1 _09180_ (.A(_04481_),
    .X(_04894_));
 sky130_fd_sc_hd__a22o_1 _09181_ (.A1(\r1.regblock[12][26] ),
    .A2(_04887_),
    .B1(_04894_),
    .B2(_04891_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_1 _09182_ (.A(_04893_),
    .X(_02101_));
 sky130_fd_sc_hd__buf_1 _09183_ (.A(_04886_),
    .X(_04895_));
 sky130_fd_sc_hd__buf_1 _09184_ (.A(_04485_),
    .X(_04896_));
 sky130_fd_sc_hd__buf_1 _09185_ (.A(_04890_),
    .X(_04897_));
 sky130_fd_sc_hd__a22o_1 _09186_ (.A1(\r1.regblock[12][25] ),
    .A2(_04895_),
    .B1(_04896_),
    .B2(_04897_),
    .X(_03126_));
 sky130_fd_sc_hd__clkbuf_1 _09187_ (.A(_04893_),
    .X(_02100_));
 sky130_fd_sc_hd__buf_1 _09188_ (.A(_04489_),
    .X(_04898_));
 sky130_fd_sc_hd__a22o_1 _09189_ (.A1(\r1.regblock[12][24] ),
    .A2(_04895_),
    .B1(_04898_),
    .B2(_04897_),
    .X(_03125_));
 sky130_fd_sc_hd__buf_1 _09190_ (.A(_04882_),
    .X(_04899_));
 sky130_fd_sc_hd__clkbuf_1 _09191_ (.A(_04899_),
    .X(_02099_));
 sky130_fd_sc_hd__buf_1 _09192_ (.A(_04493_),
    .X(_04900_));
 sky130_fd_sc_hd__a22o_1 _09193_ (.A1(\r1.regblock[12][23] ),
    .A2(_04895_),
    .B1(_04900_),
    .B2(_04897_),
    .X(_03124_));
 sky130_fd_sc_hd__clkbuf_1 _09194_ (.A(_04899_),
    .X(_02098_));
 sky130_fd_sc_hd__buf_1 _09195_ (.A(_04886_),
    .X(_04901_));
 sky130_fd_sc_hd__buf_1 _09196_ (.A(_04497_),
    .X(_04902_));
 sky130_fd_sc_hd__buf_1 _09197_ (.A(_04890_),
    .X(_04903_));
 sky130_fd_sc_hd__a22o_1 _09198_ (.A1(\r1.regblock[12][22] ),
    .A2(_04901_),
    .B1(_04902_),
    .B2(_04903_),
    .X(_03123_));
 sky130_fd_sc_hd__clkbuf_1 _09199_ (.A(_04899_),
    .X(_02097_));
 sky130_fd_sc_hd__buf_1 _09200_ (.A(_04501_),
    .X(_04904_));
 sky130_fd_sc_hd__a22o_1 _09201_ (.A1(\r1.regblock[12][21] ),
    .A2(_04901_),
    .B1(_04904_),
    .B2(_04903_),
    .X(_03122_));
 sky130_fd_sc_hd__buf_2 _09202_ (.A(_04811_),
    .X(_04905_));
 sky130_fd_sc_hd__clkbuf_2 _09203_ (.A(_04905_),
    .X(_04906_));
 sky130_fd_sc_hd__buf_1 _09204_ (.A(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__clkbuf_2 _09205_ (.A(_04907_),
    .X(_02096_));
 sky130_fd_sc_hd__buf_1 _09206_ (.A(_04505_),
    .X(_04908_));
 sky130_fd_sc_hd__a22o_1 _09207_ (.A1(\r1.regblock[12][20] ),
    .A2(_04901_),
    .B1(_04908_),
    .B2(_04903_),
    .X(_03121_));
 sky130_fd_sc_hd__clkbuf_1 _09208_ (.A(_04907_),
    .X(_02095_));
 sky130_fd_sc_hd__clkbuf_2 _09209_ (.A(_04885_),
    .X(_04909_));
 sky130_fd_sc_hd__buf_1 _09210_ (.A(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__buf_1 _09211_ (.A(_04510_),
    .X(_04911_));
 sky130_fd_sc_hd__clkbuf_2 _09212_ (.A(_04889_),
    .X(_04912_));
 sky130_fd_sc_hd__buf_1 _09213_ (.A(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__a22o_1 _09214_ (.A1(\r1.regblock[12][19] ),
    .A2(_04910_),
    .B1(_04911_),
    .B2(_04913_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_1 _09215_ (.A(_04907_),
    .X(_02094_));
 sky130_fd_sc_hd__buf_1 _09216_ (.A(_04515_),
    .X(_04914_));
 sky130_fd_sc_hd__a22o_1 _09217_ (.A1(\r1.regblock[12][18] ),
    .A2(_04910_),
    .B1(_04914_),
    .B2(_04913_),
    .X(_03119_));
 sky130_fd_sc_hd__buf_1 _09218_ (.A(_04906_),
    .X(_04915_));
 sky130_fd_sc_hd__clkbuf_1 _09219_ (.A(_04915_),
    .X(_02093_));
 sky130_fd_sc_hd__buf_1 _09220_ (.A(_04521_),
    .X(_04916_));
 sky130_fd_sc_hd__a22o_1 _09221_ (.A1(\r1.regblock[12][17] ),
    .A2(_04910_),
    .B1(_04916_),
    .B2(_04913_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_1 _09222_ (.A(_04915_),
    .X(_02092_));
 sky130_fd_sc_hd__buf_1 _09223_ (.A(_04909_),
    .X(_04917_));
 sky130_fd_sc_hd__buf_1 _09224_ (.A(_04525_),
    .X(_04918_));
 sky130_fd_sc_hd__buf_1 _09225_ (.A(_04912_),
    .X(_04919_));
 sky130_fd_sc_hd__a22o_1 _09226_ (.A1(\r1.regblock[12][16] ),
    .A2(_04917_),
    .B1(_04918_),
    .B2(_04919_),
    .X(_03117_));
 sky130_fd_sc_hd__clkbuf_1 _09227_ (.A(_04915_),
    .X(_02091_));
 sky130_fd_sc_hd__buf_1 _09228_ (.A(_04529_),
    .X(_04920_));
 sky130_fd_sc_hd__a22o_1 _09229_ (.A1(\r1.regblock[12][15] ),
    .A2(_04917_),
    .B1(_04920_),
    .B2(_04919_),
    .X(_03116_));
 sky130_fd_sc_hd__buf_1 _09230_ (.A(_04906_),
    .X(_04921_));
 sky130_fd_sc_hd__clkbuf_1 _09231_ (.A(_04921_),
    .X(_02090_));
 sky130_fd_sc_hd__buf_1 _09232_ (.A(_04533_),
    .X(_04922_));
 sky130_fd_sc_hd__a22o_1 _09233_ (.A1(\r1.regblock[12][14] ),
    .A2(_04917_),
    .B1(_04922_),
    .B2(_04919_),
    .X(_03115_));
 sky130_fd_sc_hd__clkbuf_1 _09234_ (.A(_04921_),
    .X(_02089_));
 sky130_fd_sc_hd__buf_1 _09235_ (.A(_04909_),
    .X(_04923_));
 sky130_fd_sc_hd__buf_1 _09236_ (.A(_04537_),
    .X(_04924_));
 sky130_fd_sc_hd__buf_1 _09237_ (.A(_04912_),
    .X(_04925_));
 sky130_fd_sc_hd__a22o_1 _09238_ (.A1(\r1.regblock[12][13] ),
    .A2(_04923_),
    .B1(_04924_),
    .B2(_04925_),
    .X(_03114_));
 sky130_fd_sc_hd__clkbuf_1 _09239_ (.A(_04921_),
    .X(_02088_));
 sky130_fd_sc_hd__buf_1 _09240_ (.A(_04541_),
    .X(_04926_));
 sky130_fd_sc_hd__a22o_1 _09241_ (.A1(\r1.regblock[12][12] ),
    .A2(_04923_),
    .B1(_04926_),
    .B2(_04925_),
    .X(_03113_));
 sky130_fd_sc_hd__clkbuf_2 _09242_ (.A(_04905_),
    .X(_04927_));
 sky130_fd_sc_hd__clkbuf_2 _09243_ (.A(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__clkbuf_1 _09244_ (.A(_04928_),
    .X(_02087_));
 sky130_fd_sc_hd__buf_1 _09245_ (.A(_04545_),
    .X(_04929_));
 sky130_fd_sc_hd__a22o_1 _09246_ (.A1(\r1.regblock[12][11] ),
    .A2(_04923_),
    .B1(_04929_),
    .B2(_04925_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_1 _09247_ (.A(_04928_),
    .X(_02086_));
 sky130_fd_sc_hd__buf_1 _09248_ (.A(_04885_),
    .X(_04930_));
 sky130_fd_sc_hd__buf_1 _09249_ (.A(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__buf_1 _09250_ (.A(_04550_),
    .X(_04932_));
 sky130_fd_sc_hd__buf_1 _09251_ (.A(_04889_),
    .X(_04933_));
 sky130_fd_sc_hd__buf_1 _09252_ (.A(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__a22o_1 _09253_ (.A1(\r1.regblock[12][10] ),
    .A2(_04931_),
    .B1(_04932_),
    .B2(_04934_),
    .X(_03111_));
 sky130_fd_sc_hd__clkbuf_1 _09254_ (.A(_04928_),
    .X(_02085_));
 sky130_fd_sc_hd__buf_1 _09255_ (.A(_04555_),
    .X(_04935_));
 sky130_fd_sc_hd__a22o_1 _09256_ (.A1(\r1.regblock[12][9] ),
    .A2(_04931_),
    .B1(_04935_),
    .B2(_04934_),
    .X(_03110_));
 sky130_fd_sc_hd__buf_1 _09257_ (.A(_04927_),
    .X(_04936_));
 sky130_fd_sc_hd__clkbuf_1 _09258_ (.A(_04936_),
    .X(_02084_));
 sky130_fd_sc_hd__buf_1 _09259_ (.A(_04560_),
    .X(_04937_));
 sky130_fd_sc_hd__a22o_1 _09260_ (.A1(\r1.regblock[12][8] ),
    .A2(_04931_),
    .B1(_04937_),
    .B2(_04934_),
    .X(_03109_));
 sky130_fd_sc_hd__clkbuf_1 _09261_ (.A(_04936_),
    .X(_02083_));
 sky130_fd_sc_hd__buf_1 _09262_ (.A(_04930_),
    .X(_04938_));
 sky130_fd_sc_hd__buf_1 _09263_ (.A(_04564_),
    .X(_04939_));
 sky130_fd_sc_hd__buf_1 _09264_ (.A(_04933_),
    .X(_04940_));
 sky130_fd_sc_hd__a22o_1 _09265_ (.A1(\r1.regblock[12][7] ),
    .A2(_04938_),
    .B1(_04939_),
    .B2(_04940_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _09266_ (.A(_04936_),
    .X(_02082_));
 sky130_fd_sc_hd__buf_1 _09267_ (.A(_04568_),
    .X(_04941_));
 sky130_fd_sc_hd__a22o_1 _09268_ (.A1(\r1.regblock[12][6] ),
    .A2(_04938_),
    .B1(_04941_),
    .B2(_04940_),
    .X(_03107_));
 sky130_fd_sc_hd__buf_1 _09269_ (.A(_04927_),
    .X(_04942_));
 sky130_fd_sc_hd__clkbuf_1 _09270_ (.A(_04942_),
    .X(_02081_));
 sky130_fd_sc_hd__buf_1 _09271_ (.A(_04572_),
    .X(_04943_));
 sky130_fd_sc_hd__a22o_1 _09272_ (.A1(\r1.regblock[12][5] ),
    .A2(_04938_),
    .B1(_04943_),
    .B2(_04940_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_1 _09273_ (.A(_04942_),
    .X(_02080_));
 sky130_fd_sc_hd__buf_1 _09274_ (.A(_04930_),
    .X(_04944_));
 sky130_fd_sc_hd__buf_1 _09275_ (.A(_04576_),
    .X(_04945_));
 sky130_fd_sc_hd__buf_1 _09276_ (.A(_04933_),
    .X(_04946_));
 sky130_fd_sc_hd__a22o_1 _09277_ (.A1(\r1.regblock[12][4] ),
    .A2(_04944_),
    .B1(_04945_),
    .B2(_04946_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _09278_ (.A(_04942_),
    .X(_02079_));
 sky130_fd_sc_hd__buf_1 _09279_ (.A(_04580_),
    .X(_04947_));
 sky130_fd_sc_hd__a22o_1 _09280_ (.A1(\r1.regblock[12][3] ),
    .A2(_04944_),
    .B1(_04947_),
    .B2(_04946_),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_4 _09281_ (.A(_04905_),
    .X(_04948_));
 sky130_fd_sc_hd__buf_1 _09282_ (.A(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__buf_1 _09283_ (.A(_04949_),
    .X(_02078_));
 sky130_fd_sc_hd__buf_1 _09284_ (.A(_04584_),
    .X(_04950_));
 sky130_fd_sc_hd__a22o_1 _09285_ (.A1(\r1.regblock[12][2] ),
    .A2(_04944_),
    .B1(_04950_),
    .B2(_04946_),
    .X(_03103_));
 sky130_fd_sc_hd__clkbuf_1 _09286_ (.A(_04949_),
    .X(_02077_));
 sky130_fd_sc_hd__buf_1 _09287_ (.A(_04587_),
    .X(_04951_));
 sky130_fd_sc_hd__a22o_1 _09288_ (.A1(\r1.regblock[12][1] ),
    .A2(_04875_),
    .B1(_04951_),
    .B2(_04879_),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_1 _09289_ (.A(_04949_),
    .X(_02076_));
 sky130_fd_sc_hd__buf_1 _09290_ (.A(_04590_),
    .X(_04952_));
 sky130_fd_sc_hd__a22o_1 _09291_ (.A1(\r1.regblock[12][0] ),
    .A2(_04875_),
    .B1(_04952_),
    .B2(_04879_),
    .X(_03101_));
 sky130_fd_sc_hd__buf_1 _09292_ (.A(_04948_),
    .X(_04953_));
 sky130_fd_sc_hd__clkbuf_1 _09293_ (.A(_04953_),
    .X(_02075_));
 sky130_fd_sc_hd__or3_1 _09294_ (.A(_04341_),
    .B(_04390_),
    .C(_04392_),
    .X(_04954_));
 sky130_fd_sc_hd__clkbuf_1 _09295_ (.A(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__or2_1 _09296_ (.A(_04339_),
    .B(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__buf_1 _09297_ (.A(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__buf_1 _09298_ (.A(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__inv_2 _09299_ (.A(_04956_),
    .Y(_04959_));
 sky130_fd_sc_hd__buf_1 _09300_ (.A(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__buf_1 _09301_ (.A(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__a22o_1 _09302_ (.A1(\r1.regblock[31][31] ),
    .A2(_04958_),
    .B1(_04877_),
    .B2(_04961_),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_1 _09303_ (.A(_04953_),
    .X(_02074_));
 sky130_fd_sc_hd__a22o_1 _09304_ (.A1(\r1.regblock[31][30] ),
    .A2(_04958_),
    .B1(_04881_),
    .B2(_04961_),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _09305_ (.A(_04953_),
    .X(_02073_));
 sky130_fd_sc_hd__a22o_1 _09306_ (.A1(\r1.regblock[31][29] ),
    .A2(_04958_),
    .B1(_04884_),
    .B2(_04961_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_1 _09307_ (.A(_04948_),
    .X(_04962_));
 sky130_fd_sc_hd__clkbuf_1 _09308_ (.A(_04962_),
    .X(_02072_));
 sky130_fd_sc_hd__buf_2 _09309_ (.A(_04956_),
    .X(_04963_));
 sky130_fd_sc_hd__buf_2 _09310_ (.A(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__buf_1 _09311_ (.A(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__buf_2 _09312_ (.A(_04959_),
    .X(_04966_));
 sky130_fd_sc_hd__buf_2 _09313_ (.A(_04966_),
    .X(_04967_));
 sky130_fd_sc_hd__buf_1 _09314_ (.A(_04967_),
    .X(_04968_));
 sky130_fd_sc_hd__a22o_1 _09315_ (.A1(\r1.regblock[31][28] ),
    .A2(_04965_),
    .B1(_04888_),
    .B2(_04968_),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_1 _09316_ (.A(_04962_),
    .X(_02071_));
 sky130_fd_sc_hd__a22o_1 _09317_ (.A1(\r1.regblock[31][27] ),
    .A2(_04965_),
    .B1(_04892_),
    .B2(_04968_),
    .X(_03096_));
 sky130_fd_sc_hd__clkbuf_1 _09318_ (.A(_04962_),
    .X(_02070_));
 sky130_fd_sc_hd__a22o_1 _09319_ (.A1(\r1.regblock[31][26] ),
    .A2(_04965_),
    .B1(_04894_),
    .B2(_04968_),
    .X(_03095_));
 sky130_fd_sc_hd__buf_1 _09320_ (.A(_04429_),
    .X(_04969_));
 sky130_fd_sc_hd__clkbuf_1 _09321_ (.A(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__buf_1 _09322_ (.A(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__clkbuf_4 _09323_ (.A(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__buf_1 _09324_ (.A(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__clkbuf_1 _09325_ (.A(_04973_),
    .X(_02069_));
 sky130_fd_sc_hd__buf_1 _09326_ (.A(_04964_),
    .X(_04974_));
 sky130_fd_sc_hd__buf_1 _09327_ (.A(_04967_),
    .X(_04975_));
 sky130_fd_sc_hd__a22o_1 _09328_ (.A1(\r1.regblock[31][25] ),
    .A2(_04974_),
    .B1(_04896_),
    .B2(_04975_),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_1 _09329_ (.A(_04973_),
    .X(_02068_));
 sky130_fd_sc_hd__a22o_1 _09330_ (.A1(\r1.regblock[31][24] ),
    .A2(_04974_),
    .B1(_04898_),
    .B2(_04975_),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_1 _09331_ (.A(_04973_),
    .X(_02067_));
 sky130_fd_sc_hd__a22o_1 _09332_ (.A1(\r1.regblock[31][23] ),
    .A2(_04974_),
    .B1(_04900_),
    .B2(_04975_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_1 _09333_ (.A(_04972_),
    .X(_04976_));
 sky130_fd_sc_hd__clkbuf_1 _09334_ (.A(_04976_),
    .X(_02066_));
 sky130_fd_sc_hd__buf_1 _09335_ (.A(_04964_),
    .X(_04977_));
 sky130_fd_sc_hd__buf_1 _09336_ (.A(_04967_),
    .X(_04978_));
 sky130_fd_sc_hd__a22o_1 _09337_ (.A1(\r1.regblock[31][22] ),
    .A2(_04977_),
    .B1(_04902_),
    .B2(_04978_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_1 _09338_ (.A(_04976_),
    .X(_02065_));
 sky130_fd_sc_hd__a22o_1 _09339_ (.A1(\r1.regblock[31][21] ),
    .A2(_04977_),
    .B1(_04904_),
    .B2(_04978_),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _09340_ (.A(_04976_),
    .X(_02064_));
 sky130_fd_sc_hd__a22o_1 _09341_ (.A1(\r1.regblock[31][20] ),
    .A2(_04977_),
    .B1(_04908_),
    .B2(_04978_),
    .X(_03089_));
 sky130_fd_sc_hd__buf_1 _09342_ (.A(_04972_),
    .X(_04979_));
 sky130_fd_sc_hd__clkbuf_1 _09343_ (.A(_04979_),
    .X(_02063_));
 sky130_fd_sc_hd__buf_2 _09344_ (.A(_04963_),
    .X(_04980_));
 sky130_fd_sc_hd__buf_1 _09345_ (.A(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__buf_2 _09346_ (.A(_04966_),
    .X(_04982_));
 sky130_fd_sc_hd__buf_1 _09347_ (.A(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__a22o_1 _09348_ (.A1(\r1.regblock[31][19] ),
    .A2(_04981_),
    .B1(_04911_),
    .B2(_04983_),
    .X(_03088_));
 sky130_fd_sc_hd__clkbuf_1 _09349_ (.A(_04979_),
    .X(_02062_));
 sky130_fd_sc_hd__a22o_1 _09350_ (.A1(\r1.regblock[31][18] ),
    .A2(_04981_),
    .B1(_04914_),
    .B2(_04983_),
    .X(_03087_));
 sky130_fd_sc_hd__clkbuf_1 _09351_ (.A(_04979_),
    .X(_02061_));
 sky130_fd_sc_hd__a22o_1 _09352_ (.A1(\r1.regblock[31][17] ),
    .A2(_04981_),
    .B1(_04916_),
    .B2(_04983_),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_4 _09353_ (.A(_04971_),
    .X(_04984_));
 sky130_fd_sc_hd__buf_1 _09354_ (.A(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__clkbuf_1 _09355_ (.A(_04985_),
    .X(_02060_));
 sky130_fd_sc_hd__buf_1 _09356_ (.A(_04980_),
    .X(_04986_));
 sky130_fd_sc_hd__buf_1 _09357_ (.A(_04982_),
    .X(_04987_));
 sky130_fd_sc_hd__a22o_1 _09358_ (.A1(\r1.regblock[31][16] ),
    .A2(_04986_),
    .B1(_04918_),
    .B2(_04987_),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_1 _09359_ (.A(_04985_),
    .X(_02059_));
 sky130_fd_sc_hd__a22o_1 _09360_ (.A1(\r1.regblock[31][15] ),
    .A2(_04986_),
    .B1(_04920_),
    .B2(_04987_),
    .X(_03084_));
 sky130_fd_sc_hd__clkbuf_1 _09361_ (.A(_04985_),
    .X(_02058_));
 sky130_fd_sc_hd__a22o_1 _09362_ (.A1(\r1.regblock[31][14] ),
    .A2(_04986_),
    .B1(_04922_),
    .B2(_04987_),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_1 _09363_ (.A(_04984_),
    .X(_04988_));
 sky130_fd_sc_hd__clkbuf_1 _09364_ (.A(_04988_),
    .X(_02057_));
 sky130_fd_sc_hd__buf_1 _09365_ (.A(_04980_),
    .X(_04989_));
 sky130_fd_sc_hd__buf_1 _09366_ (.A(_04982_),
    .X(_04990_));
 sky130_fd_sc_hd__a22o_1 _09367_ (.A1(\r1.regblock[31][13] ),
    .A2(_04989_),
    .B1(_04924_),
    .B2(_04990_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _09368_ (.A(_04988_),
    .X(_02056_));
 sky130_fd_sc_hd__a22o_1 _09369_ (.A1(\r1.regblock[31][12] ),
    .A2(_04989_),
    .B1(_04926_),
    .B2(_04990_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_1 _09370_ (.A(_04988_),
    .X(_02055_));
 sky130_fd_sc_hd__a22o_1 _09371_ (.A1(\r1.regblock[31][11] ),
    .A2(_04989_),
    .B1(_04929_),
    .B2(_04990_),
    .X(_03080_));
 sky130_fd_sc_hd__buf_1 _09372_ (.A(_04984_),
    .X(_04991_));
 sky130_fd_sc_hd__clkbuf_1 _09373_ (.A(_04991_),
    .X(_02054_));
 sky130_fd_sc_hd__clkbuf_2 _09374_ (.A(_04963_),
    .X(_04992_));
 sky130_fd_sc_hd__buf_1 _09375_ (.A(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__clkbuf_2 _09376_ (.A(_04966_),
    .X(_04994_));
 sky130_fd_sc_hd__buf_1 _09377_ (.A(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__a22o_1 _09378_ (.A1(\r1.regblock[31][10] ),
    .A2(_04993_),
    .B1(_04932_),
    .B2(_04995_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _09379_ (.A(_04991_),
    .X(_02053_));
 sky130_fd_sc_hd__a22o_1 _09380_ (.A1(\r1.regblock[31][9] ),
    .A2(_04993_),
    .B1(_04935_),
    .B2(_04995_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_1 _09381_ (.A(_04991_),
    .X(_02052_));
 sky130_fd_sc_hd__a22o_1 _09382_ (.A1(\r1.regblock[31][8] ),
    .A2(_04993_),
    .B1(_04937_),
    .B2(_04995_),
    .X(_03077_));
 sky130_fd_sc_hd__clkbuf_2 _09383_ (.A(_04971_),
    .X(_04996_));
 sky130_fd_sc_hd__buf_1 _09384_ (.A(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__clkbuf_1 _09385_ (.A(_04997_),
    .X(_02051_));
 sky130_fd_sc_hd__buf_1 _09386_ (.A(_04992_),
    .X(_04998_));
 sky130_fd_sc_hd__buf_1 _09387_ (.A(_04994_),
    .X(_04999_));
 sky130_fd_sc_hd__a22o_1 _09388_ (.A1(\r1.regblock[31][7] ),
    .A2(_04998_),
    .B1(_04939_),
    .B2(_04999_),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_1 _09389_ (.A(_04997_),
    .X(_02050_));
 sky130_fd_sc_hd__a22o_1 _09390_ (.A1(\r1.regblock[31][6] ),
    .A2(_04998_),
    .B1(_04941_),
    .B2(_04999_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_1 _09391_ (.A(_04997_),
    .X(_02049_));
 sky130_fd_sc_hd__a22o_1 _09392_ (.A1(\r1.regblock[31][5] ),
    .A2(_04998_),
    .B1(_04943_),
    .B2(_04999_),
    .X(_03074_));
 sky130_fd_sc_hd__buf_1 _09393_ (.A(_04996_),
    .X(_05000_));
 sky130_fd_sc_hd__clkbuf_1 _09394_ (.A(_05000_),
    .X(_02048_));
 sky130_fd_sc_hd__buf_1 _09395_ (.A(_04992_),
    .X(_05001_));
 sky130_fd_sc_hd__buf_1 _09396_ (.A(_04994_),
    .X(_05002_));
 sky130_fd_sc_hd__a22o_1 _09397_ (.A1(\r1.regblock[31][4] ),
    .A2(_05001_),
    .B1(_04945_),
    .B2(_05002_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_1 _09398_ (.A(_05000_),
    .X(_02047_));
 sky130_fd_sc_hd__a22o_1 _09399_ (.A1(\r1.regblock[31][3] ),
    .A2(_05001_),
    .B1(_04947_),
    .B2(_05002_),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_1 _09400_ (.A(_05000_),
    .X(_02046_));
 sky130_fd_sc_hd__a22o_1 _09401_ (.A1(\r1.regblock[31][2] ),
    .A2(_05001_),
    .B1(_04950_),
    .B2(_05002_),
    .X(_03071_));
 sky130_fd_sc_hd__buf_1 _09402_ (.A(_04996_),
    .X(_05003_));
 sky130_fd_sc_hd__clkbuf_1 _09403_ (.A(_05003_),
    .X(_02045_));
 sky130_fd_sc_hd__a22o_1 _09404_ (.A1(\r1.regblock[31][1] ),
    .A2(_04957_),
    .B1(_04951_),
    .B2(_04960_),
    .X(_03070_));
 sky130_fd_sc_hd__clkbuf_1 _09405_ (.A(_05003_),
    .X(_02044_));
 sky130_fd_sc_hd__a22o_1 _09406_ (.A1(\r1.regblock[31][0] ),
    .A2(_04957_),
    .B1(_04952_),
    .B2(_04960_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _09407_ (.A(_05003_),
    .X(_02043_));
 sky130_fd_sc_hd__or2_1 _09408_ (.A(_04641_),
    .B(_04955_),
    .X(_05004_));
 sky130_fd_sc_hd__buf_1 _09409_ (.A(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__buf_1 _09410_ (.A(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__inv_2 _09411_ (.A(_05004_),
    .Y(_05007_));
 sky130_fd_sc_hd__buf_1 _09412_ (.A(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__buf_1 _09413_ (.A(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__a22o_1 _09414_ (.A1(\r1.regblock[29][31] ),
    .A2(_05006_),
    .B1(_04877_),
    .B2(_05009_),
    .X(_03068_));
 sky130_fd_sc_hd__buf_1 _09415_ (.A(_04970_),
    .X(_05010_));
 sky130_fd_sc_hd__buf_2 _09416_ (.A(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__clkbuf_2 _09417_ (.A(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__clkbuf_1 _09418_ (.A(_05012_),
    .X(_02042_));
 sky130_fd_sc_hd__a22o_1 _09419_ (.A1(\r1.regblock[29][30] ),
    .A2(_05006_),
    .B1(_04881_),
    .B2(_05009_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_1 _09420_ (.A(_05012_),
    .X(_02041_));
 sky130_fd_sc_hd__a22o_1 _09421_ (.A1(\r1.regblock[29][29] ),
    .A2(_05006_),
    .B1(_04884_),
    .B2(_05009_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_1 _09422_ (.A(_05012_),
    .X(_02040_));
 sky130_fd_sc_hd__buf_2 _09423_ (.A(_05004_),
    .X(_05013_));
 sky130_fd_sc_hd__clkbuf_2 _09424_ (.A(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__buf_1 _09425_ (.A(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__buf_2 _09426_ (.A(_05007_),
    .X(_05016_));
 sky130_fd_sc_hd__clkbuf_2 _09427_ (.A(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__buf_1 _09428_ (.A(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__a22o_1 _09429_ (.A1(\r1.regblock[29][28] ),
    .A2(_05015_),
    .B1(_04888_),
    .B2(_05018_),
    .X(_03065_));
 sky130_fd_sc_hd__buf_1 _09430_ (.A(_05011_),
    .X(_05019_));
 sky130_fd_sc_hd__clkbuf_1 _09431_ (.A(_05019_),
    .X(_02039_));
 sky130_fd_sc_hd__a22o_1 _09432_ (.A1(\r1.regblock[29][27] ),
    .A2(_05015_),
    .B1(_04892_),
    .B2(_05018_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _09433_ (.A(_05019_),
    .X(_02038_));
 sky130_fd_sc_hd__a22o_1 _09434_ (.A1(\r1.regblock[29][26] ),
    .A2(_05015_),
    .B1(_04894_),
    .B2(_05018_),
    .X(_03063_));
 sky130_fd_sc_hd__clkbuf_1 _09435_ (.A(_05019_),
    .X(_02037_));
 sky130_fd_sc_hd__buf_1 _09436_ (.A(_05014_),
    .X(_05020_));
 sky130_fd_sc_hd__buf_1 _09437_ (.A(_05017_),
    .X(_05021_));
 sky130_fd_sc_hd__a22o_1 _09438_ (.A1(\r1.regblock[29][25] ),
    .A2(_05020_),
    .B1(_04896_),
    .B2(_05021_),
    .X(_03062_));
 sky130_fd_sc_hd__buf_1 _09439_ (.A(_05011_),
    .X(_05022_));
 sky130_fd_sc_hd__clkbuf_1 _09440_ (.A(_05022_),
    .X(_02036_));
 sky130_fd_sc_hd__a22o_1 _09441_ (.A1(\r1.regblock[29][24] ),
    .A2(_05020_),
    .B1(_04898_),
    .B2(_05021_),
    .X(_03061_));
 sky130_fd_sc_hd__clkbuf_1 _09442_ (.A(_05022_),
    .X(_02035_));
 sky130_fd_sc_hd__a22o_1 _09443_ (.A1(\r1.regblock[29][23] ),
    .A2(_05020_),
    .B1(_04900_),
    .B2(_05021_),
    .X(_03060_));
 sky130_fd_sc_hd__clkbuf_1 _09444_ (.A(_05022_),
    .X(_02034_));
 sky130_fd_sc_hd__buf_1 _09445_ (.A(_05014_),
    .X(_05023_));
 sky130_fd_sc_hd__buf_1 _09446_ (.A(_05017_),
    .X(_05024_));
 sky130_fd_sc_hd__a22o_1 _09447_ (.A1(\r1.regblock[29][22] ),
    .A2(_05023_),
    .B1(_04902_),
    .B2(_05024_),
    .X(_03059_));
 sky130_fd_sc_hd__buf_2 _09448_ (.A(_05010_),
    .X(_05025_));
 sky130_fd_sc_hd__buf_2 _09449_ (.A(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__clkbuf_1 _09450_ (.A(_05026_),
    .X(_02033_));
 sky130_fd_sc_hd__a22o_1 _09451_ (.A1(\r1.regblock[29][21] ),
    .A2(_05023_),
    .B1(_04904_),
    .B2(_05024_),
    .X(_03058_));
 sky130_fd_sc_hd__clkbuf_1 _09452_ (.A(_05026_),
    .X(_02032_));
 sky130_fd_sc_hd__a22o_1 _09453_ (.A1(\r1.regblock[29][20] ),
    .A2(_05023_),
    .B1(_04908_),
    .B2(_05024_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_1 _09454_ (.A(_05026_),
    .X(_02031_));
 sky130_fd_sc_hd__buf_2 _09455_ (.A(_05013_),
    .X(_05027_));
 sky130_fd_sc_hd__buf_1 _09456_ (.A(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__buf_2 _09457_ (.A(_05016_),
    .X(_05029_));
 sky130_fd_sc_hd__buf_1 _09458_ (.A(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__a22o_1 _09459_ (.A1(\r1.regblock[29][19] ),
    .A2(_05028_),
    .B1(_04911_),
    .B2(_05030_),
    .X(_03056_));
 sky130_fd_sc_hd__buf_1 _09460_ (.A(_05025_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_1 _09461_ (.A(_05031_),
    .X(_02030_));
 sky130_fd_sc_hd__a22o_1 _09462_ (.A1(\r1.regblock[29][18] ),
    .A2(_05028_),
    .B1(_04914_),
    .B2(_05030_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_1 _09463_ (.A(_05031_),
    .X(_02029_));
 sky130_fd_sc_hd__a22o_1 _09464_ (.A1(\r1.regblock[29][17] ),
    .A2(_05028_),
    .B1(_04916_),
    .B2(_05030_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _09465_ (.A(_05031_),
    .X(_02028_));
 sky130_fd_sc_hd__buf_1 _09466_ (.A(_05027_),
    .X(_05032_));
 sky130_fd_sc_hd__buf_1 _09467_ (.A(_05029_),
    .X(_05033_));
 sky130_fd_sc_hd__a22o_1 _09468_ (.A1(\r1.regblock[29][16] ),
    .A2(_05032_),
    .B1(_04918_),
    .B2(_05033_),
    .X(_03053_));
 sky130_fd_sc_hd__buf_1 _09469_ (.A(_05025_),
    .X(_05034_));
 sky130_fd_sc_hd__clkbuf_1 _09470_ (.A(_05034_),
    .X(_02027_));
 sky130_fd_sc_hd__a22o_1 _09471_ (.A1(\r1.regblock[29][15] ),
    .A2(_05032_),
    .B1(_04920_),
    .B2(_05033_),
    .X(_03052_));
 sky130_fd_sc_hd__clkbuf_1 _09472_ (.A(_05034_),
    .X(_02026_));
 sky130_fd_sc_hd__a22o_1 _09473_ (.A1(\r1.regblock[29][14] ),
    .A2(_05032_),
    .B1(_04922_),
    .B2(_05033_),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_1 _09474_ (.A(_05034_),
    .X(_02025_));
 sky130_fd_sc_hd__buf_1 _09475_ (.A(_05027_),
    .X(_05035_));
 sky130_fd_sc_hd__buf_1 _09476_ (.A(_05029_),
    .X(_05036_));
 sky130_fd_sc_hd__a22o_1 _09477_ (.A1(\r1.regblock[29][13] ),
    .A2(_05035_),
    .B1(_04924_),
    .B2(_05036_),
    .X(_03050_));
 sky130_fd_sc_hd__buf_1 _09478_ (.A(_05010_),
    .X(_05037_));
 sky130_fd_sc_hd__buf_2 _09479_ (.A(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__clkbuf_1 _09480_ (.A(_05038_),
    .X(_02024_));
 sky130_fd_sc_hd__a22o_1 _09481_ (.A1(\r1.regblock[29][12] ),
    .A2(_05035_),
    .B1(_04926_),
    .B2(_05036_),
    .X(_03049_));
 sky130_fd_sc_hd__clkbuf_1 _09482_ (.A(_05038_),
    .X(_02023_));
 sky130_fd_sc_hd__a22o_1 _09483_ (.A1(\r1.regblock[29][11] ),
    .A2(_05035_),
    .B1(_04929_),
    .B2(_05036_),
    .X(_03048_));
 sky130_fd_sc_hd__clkbuf_1 _09484_ (.A(_05038_),
    .X(_02022_));
 sky130_fd_sc_hd__buf_1 _09485_ (.A(_05013_),
    .X(_05039_));
 sky130_fd_sc_hd__buf_1 _09486_ (.A(_05039_),
    .X(_05040_));
 sky130_fd_sc_hd__buf_1 _09487_ (.A(_05016_),
    .X(_05041_));
 sky130_fd_sc_hd__buf_1 _09488_ (.A(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__a22o_1 _09489_ (.A1(\r1.regblock[29][10] ),
    .A2(_05040_),
    .B1(_04932_),
    .B2(_05042_),
    .X(_03047_));
 sky130_fd_sc_hd__buf_1 _09490_ (.A(_05037_),
    .X(_05043_));
 sky130_fd_sc_hd__clkbuf_1 _09491_ (.A(_05043_),
    .X(_02021_));
 sky130_fd_sc_hd__a22o_1 _09492_ (.A1(\r1.regblock[29][9] ),
    .A2(_05040_),
    .B1(_04935_),
    .B2(_05042_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_1 _09493_ (.A(_05043_),
    .X(_02020_));
 sky130_fd_sc_hd__a22o_1 _09494_ (.A1(\r1.regblock[29][8] ),
    .A2(_05040_),
    .B1(_04937_),
    .B2(_05042_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_1 _09495_ (.A(_05043_),
    .X(_02019_));
 sky130_fd_sc_hd__buf_1 _09496_ (.A(_05039_),
    .X(_05044_));
 sky130_fd_sc_hd__buf_1 _09497_ (.A(_05041_),
    .X(_05045_));
 sky130_fd_sc_hd__a22o_1 _09498_ (.A1(\r1.regblock[29][7] ),
    .A2(_05044_),
    .B1(_04939_),
    .B2(_05045_),
    .X(_03044_));
 sky130_fd_sc_hd__buf_1 _09499_ (.A(_05037_),
    .X(_05046_));
 sky130_fd_sc_hd__clkbuf_1 _09500_ (.A(_05046_),
    .X(_02018_));
 sky130_fd_sc_hd__a22o_1 _09501_ (.A1(\r1.regblock[29][6] ),
    .A2(_05044_),
    .B1(_04941_),
    .B2(_05045_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _09502_ (.A(_05046_),
    .X(_02017_));
 sky130_fd_sc_hd__a22o_1 _09503_ (.A1(\r1.regblock[29][5] ),
    .A2(_05044_),
    .B1(_04943_),
    .B2(_05045_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _09504_ (.A(_05046_),
    .X(_02016_));
 sky130_fd_sc_hd__buf_1 _09505_ (.A(_05039_),
    .X(_05047_));
 sky130_fd_sc_hd__buf_1 _09506_ (.A(_05041_),
    .X(_05048_));
 sky130_fd_sc_hd__a22o_1 _09507_ (.A1(\r1.regblock[29][4] ),
    .A2(_05047_),
    .B1(_04945_),
    .B2(_05048_),
    .X(_03041_));
 sky130_fd_sc_hd__buf_2 _09508_ (.A(_04970_),
    .X(_05049_));
 sky130_fd_sc_hd__clkbuf_2 _09509_ (.A(_05049_),
    .X(_05050_));
 sky130_fd_sc_hd__clkbuf_2 _09510_ (.A(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__clkbuf_1 _09511_ (.A(_05051_),
    .X(_02015_));
 sky130_fd_sc_hd__a22o_1 _09512_ (.A1(\r1.regblock[29][3] ),
    .A2(_05047_),
    .B1(_04947_),
    .B2(_05048_),
    .X(_03040_));
 sky130_fd_sc_hd__clkbuf_1 _09513_ (.A(_05051_),
    .X(_02014_));
 sky130_fd_sc_hd__a22o_1 _09514_ (.A1(\r1.regblock[29][2] ),
    .A2(_05047_),
    .B1(_04950_),
    .B2(_05048_),
    .X(_03039_));
 sky130_fd_sc_hd__clkbuf_1 _09515_ (.A(_05051_),
    .X(_02013_));
 sky130_fd_sc_hd__a22o_1 _09516_ (.A1(\r1.regblock[29][1] ),
    .A2(_05005_),
    .B1(_04951_),
    .B2(_05008_),
    .X(_03038_));
 sky130_fd_sc_hd__buf_1 _09517_ (.A(_05050_),
    .X(_05052_));
 sky130_fd_sc_hd__clkbuf_1 _09518_ (.A(_05052_),
    .X(_02012_));
 sky130_fd_sc_hd__a22o_1 _09519_ (.A1(\r1.regblock[29][0] ),
    .A2(_05005_),
    .B1(_04952_),
    .B2(_05008_),
    .X(_03037_));
 sky130_fd_sc_hd__clkbuf_1 _09520_ (.A(_05052_),
    .X(_02011_));
 sky130_fd_sc_hd__buf_1 _09521_ (.A(_04448_),
    .X(_05053_));
 sky130_fd_sc_hd__buf_1 _09522_ (.A(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__or2_1 _09523_ (.A(_05054_),
    .B(_04955_),
    .X(_05055_));
 sky130_fd_sc_hd__buf_1 _09524_ (.A(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__buf_1 _09525_ (.A(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__buf_1 _09526_ (.A(_04453_),
    .X(_05058_));
 sky130_fd_sc_hd__buf_1 _09527_ (.A(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__inv_2 _09528_ (.A(_05055_),
    .Y(_05060_));
 sky130_fd_sc_hd__buf_1 _09529_ (.A(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__buf_1 _09530_ (.A(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__a22o_1 _09531_ (.A1(\r1.regblock[30][31] ),
    .A2(_05057_),
    .B1(_05059_),
    .B2(_05062_),
    .X(_03036_));
 sky130_fd_sc_hd__clkbuf_1 _09532_ (.A(_05052_),
    .X(_02010_));
 sky130_fd_sc_hd__buf_1 _09533_ (.A(_04459_),
    .X(_05063_));
 sky130_fd_sc_hd__buf_1 _09534_ (.A(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__a22o_1 _09535_ (.A1(\r1.regblock[30][30] ),
    .A2(_05057_),
    .B1(_05064_),
    .B2(_05062_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_2 _09536_ (.A(_05050_),
    .X(_05065_));
 sky130_fd_sc_hd__clkbuf_1 _09537_ (.A(_05065_),
    .X(_02009_));
 sky130_fd_sc_hd__buf_1 _09538_ (.A(_04463_),
    .X(_05066_));
 sky130_fd_sc_hd__buf_1 _09539_ (.A(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__a22o_1 _09540_ (.A1(\r1.regblock[30][29] ),
    .A2(_05057_),
    .B1(_05067_),
    .B2(_05062_),
    .X(_03034_));
 sky130_fd_sc_hd__clkbuf_1 _09541_ (.A(_05065_),
    .X(_02008_));
 sky130_fd_sc_hd__buf_2 _09542_ (.A(_05055_),
    .X(_05068_));
 sky130_fd_sc_hd__buf_2 _09543_ (.A(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__buf_1 _09544_ (.A(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__buf_1 _09545_ (.A(_04469_),
    .X(_05071_));
 sky130_fd_sc_hd__buf_1 _09546_ (.A(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__buf_2 _09547_ (.A(_05060_),
    .X(_05073_));
 sky130_fd_sc_hd__buf_2 _09548_ (.A(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__buf_1 _09549_ (.A(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__a22o_1 _09550_ (.A1(\r1.regblock[30][28] ),
    .A2(_05070_),
    .B1(_05072_),
    .B2(_05075_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_1 _09551_ (.A(_05065_),
    .X(_02007_));
 sky130_fd_sc_hd__buf_1 _09552_ (.A(_04475_),
    .X(_05076_));
 sky130_fd_sc_hd__buf_1 _09553_ (.A(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__a22o_1 _09554_ (.A1(\r1.regblock[30][27] ),
    .A2(_05070_),
    .B1(_05077_),
    .B2(_05075_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_2 _09555_ (.A(_05049_),
    .X(_05078_));
 sky130_fd_sc_hd__clkbuf_2 _09556_ (.A(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__clkbuf_1 _09557_ (.A(_05079_),
    .X(_02006_));
 sky130_fd_sc_hd__buf_1 _09558_ (.A(_04480_),
    .X(_05080_));
 sky130_fd_sc_hd__buf_1 _09559_ (.A(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__a22o_1 _09560_ (.A1(\r1.regblock[30][26] ),
    .A2(_05070_),
    .B1(_05081_),
    .B2(_05075_),
    .X(_03031_));
 sky130_fd_sc_hd__clkbuf_1 _09561_ (.A(_05079_),
    .X(_02005_));
 sky130_fd_sc_hd__buf_1 _09562_ (.A(_05069_),
    .X(_05082_));
 sky130_fd_sc_hd__buf_1 _09563_ (.A(_04484_),
    .X(_05083_));
 sky130_fd_sc_hd__buf_1 _09564_ (.A(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__buf_1 _09565_ (.A(_05074_),
    .X(_05085_));
 sky130_fd_sc_hd__a22o_1 _09566_ (.A1(\r1.regblock[30][25] ),
    .A2(_05082_),
    .B1(_05084_),
    .B2(_05085_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _09567_ (.A(_05079_),
    .X(_02004_));
 sky130_fd_sc_hd__buf_1 _09568_ (.A(_04488_),
    .X(_05086_));
 sky130_fd_sc_hd__buf_1 _09569_ (.A(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__a22o_1 _09570_ (.A1(\r1.regblock[30][24] ),
    .A2(_05082_),
    .B1(_05087_),
    .B2(_05085_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_2 _09571_ (.A(_05078_),
    .X(_05088_));
 sky130_fd_sc_hd__clkbuf_1 _09572_ (.A(_05088_),
    .X(_02003_));
 sky130_fd_sc_hd__buf_1 _09573_ (.A(_04492_),
    .X(_05089_));
 sky130_fd_sc_hd__buf_1 _09574_ (.A(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__a22o_1 _09575_ (.A1(\r1.regblock[30][23] ),
    .A2(_05082_),
    .B1(_05090_),
    .B2(_05085_),
    .X(_03028_));
 sky130_fd_sc_hd__clkbuf_1 _09576_ (.A(_05088_),
    .X(_02002_));
 sky130_fd_sc_hd__buf_1 _09577_ (.A(_05069_),
    .X(_05091_));
 sky130_fd_sc_hd__buf_1 _09578_ (.A(_04496_),
    .X(_05092_));
 sky130_fd_sc_hd__buf_1 _09579_ (.A(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__buf_1 _09580_ (.A(_05074_),
    .X(_05094_));
 sky130_fd_sc_hd__a22o_1 _09581_ (.A1(\r1.regblock[30][22] ),
    .A2(_05091_),
    .B1(_05093_),
    .B2(_05094_),
    .X(_03027_));
 sky130_fd_sc_hd__clkbuf_1 _09582_ (.A(_05088_),
    .X(_02001_));
 sky130_fd_sc_hd__buf_1 _09583_ (.A(_04500_),
    .X(_05095_));
 sky130_fd_sc_hd__buf_1 _09584_ (.A(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__a22o_1 _09585_ (.A1(\r1.regblock[30][21] ),
    .A2(_05091_),
    .B1(_05096_),
    .B2(_05094_),
    .X(_03026_));
 sky130_fd_sc_hd__buf_2 _09586_ (.A(_05078_),
    .X(_05097_));
 sky130_fd_sc_hd__clkbuf_1 _09587_ (.A(_05097_),
    .X(_02000_));
 sky130_fd_sc_hd__buf_1 _09588_ (.A(_04504_),
    .X(_05098_));
 sky130_fd_sc_hd__buf_1 _09589_ (.A(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__a22o_1 _09590_ (.A1(\r1.regblock[30][20] ),
    .A2(_05091_),
    .B1(_05099_),
    .B2(_05094_),
    .X(_03025_));
 sky130_fd_sc_hd__clkbuf_1 _09591_ (.A(_05097_),
    .X(_01999_));
 sky130_fd_sc_hd__buf_2 _09592_ (.A(_05068_),
    .X(_05100_));
 sky130_fd_sc_hd__buf_1 _09593_ (.A(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__buf_1 _09594_ (.A(_04509_),
    .X(_05102_));
 sky130_fd_sc_hd__buf_1 _09595_ (.A(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__buf_2 _09596_ (.A(_05073_),
    .X(_05104_));
 sky130_fd_sc_hd__buf_1 _09597_ (.A(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__a22o_1 _09598_ (.A1(\r1.regblock[30][19] ),
    .A2(_05101_),
    .B1(_05103_),
    .B2(_05105_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_1 _09599_ (.A(_05097_),
    .X(_01998_));
 sky130_fd_sc_hd__buf_1 _09600_ (.A(_04514_),
    .X(_05106_));
 sky130_fd_sc_hd__buf_1 _09601_ (.A(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__a22o_1 _09602_ (.A1(\r1.regblock[30][18] ),
    .A2(_05101_),
    .B1(_05107_),
    .B2(_05105_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_4 _09603_ (.A(_05049_),
    .X(_05108_));
 sky130_fd_sc_hd__buf_1 _09604_ (.A(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__clkbuf_1 _09605_ (.A(_05109_),
    .X(_01997_));
 sky130_fd_sc_hd__buf_1 _09606_ (.A(_04520_),
    .X(_05110_));
 sky130_fd_sc_hd__buf_1 _09607_ (.A(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__a22o_1 _09608_ (.A1(\r1.regblock[30][17] ),
    .A2(_05101_),
    .B1(_05111_),
    .B2(_05105_),
    .X(_03022_));
 sky130_fd_sc_hd__clkbuf_1 _09609_ (.A(_05109_),
    .X(_01996_));
 sky130_fd_sc_hd__buf_1 _09610_ (.A(_05100_),
    .X(_05112_));
 sky130_fd_sc_hd__buf_1 _09611_ (.A(_04524_),
    .X(_05113_));
 sky130_fd_sc_hd__buf_1 _09612_ (.A(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__buf_1 _09613_ (.A(_05104_),
    .X(_05115_));
 sky130_fd_sc_hd__a22o_1 _09614_ (.A1(\r1.regblock[30][16] ),
    .A2(_05112_),
    .B1(_05114_),
    .B2(_05115_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_1 _09615_ (.A(_05109_),
    .X(_01995_));
 sky130_fd_sc_hd__buf_1 _09616_ (.A(_04528_),
    .X(_05116_));
 sky130_fd_sc_hd__buf_1 _09617_ (.A(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__a22o_1 _09618_ (.A1(\r1.regblock[30][15] ),
    .A2(_05112_),
    .B1(_05117_),
    .B2(_05115_),
    .X(_03020_));
 sky130_fd_sc_hd__buf_1 _09619_ (.A(_05108_),
    .X(_05118_));
 sky130_fd_sc_hd__clkbuf_1 _09620_ (.A(_05118_),
    .X(_01994_));
 sky130_fd_sc_hd__buf_1 _09621_ (.A(_04532_),
    .X(_05119_));
 sky130_fd_sc_hd__buf_1 _09622_ (.A(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__a22o_1 _09623_ (.A1(\r1.regblock[30][14] ),
    .A2(_05112_),
    .B1(_05120_),
    .B2(_05115_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_1 _09624_ (.A(_05118_),
    .X(_01993_));
 sky130_fd_sc_hd__buf_1 _09625_ (.A(_05100_),
    .X(_05121_));
 sky130_fd_sc_hd__buf_1 _09626_ (.A(_04536_),
    .X(_05122_));
 sky130_fd_sc_hd__buf_1 _09627_ (.A(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__buf_1 _09628_ (.A(_05104_),
    .X(_05124_));
 sky130_fd_sc_hd__a22o_1 _09629_ (.A1(\r1.regblock[30][13] ),
    .A2(_05121_),
    .B1(_05123_),
    .B2(_05124_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_1 _09630_ (.A(_05118_),
    .X(_01992_));
 sky130_fd_sc_hd__buf_1 _09631_ (.A(_04540_),
    .X(_05125_));
 sky130_fd_sc_hd__buf_1 _09632_ (.A(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__a22o_1 _09633_ (.A1(\r1.regblock[30][12] ),
    .A2(_05121_),
    .B1(_05126_),
    .B2(_05124_),
    .X(_03017_));
 sky130_fd_sc_hd__buf_1 _09634_ (.A(_05108_),
    .X(_05127_));
 sky130_fd_sc_hd__buf_1 _09635_ (.A(_05127_),
    .X(_01991_));
 sky130_fd_sc_hd__buf_1 _09636_ (.A(_04544_),
    .X(_05128_));
 sky130_fd_sc_hd__buf_1 _09637_ (.A(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__a22o_1 _09638_ (.A1(\r1.regblock[30][11] ),
    .A2(_05121_),
    .B1(_05129_),
    .B2(_05124_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_1 _09639_ (.A(_05127_),
    .X(_01990_));
 sky130_fd_sc_hd__buf_1 _09640_ (.A(_05068_),
    .X(_05130_));
 sky130_fd_sc_hd__buf_1 _09641_ (.A(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__buf_1 _09642_ (.A(_04549_),
    .X(_05132_));
 sky130_fd_sc_hd__buf_1 _09643_ (.A(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__buf_1 _09644_ (.A(_05073_),
    .X(_05134_));
 sky130_fd_sc_hd__buf_1 _09645_ (.A(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__a22o_1 _09646_ (.A1(\r1.regblock[30][10] ),
    .A2(_05131_),
    .B1(_05133_),
    .B2(_05135_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_1 _09647_ (.A(_05127_),
    .X(_01989_));
 sky130_fd_sc_hd__buf_1 _09648_ (.A(_04554_),
    .X(_05136_));
 sky130_fd_sc_hd__buf_1 _09649_ (.A(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__a22o_1 _09650_ (.A1(\r1.regblock[30][9] ),
    .A2(_05131_),
    .B1(_05137_),
    .B2(_05135_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_1 _09651_ (.A(_04969_),
    .X(_05138_));
 sky130_fd_sc_hd__buf_1 _09652_ (.A(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__clkbuf_2 _09653_ (.A(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__buf_1 _09654_ (.A(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__clkbuf_1 _09655_ (.A(_05141_),
    .X(_01988_));
 sky130_fd_sc_hd__buf_1 _09656_ (.A(_04559_),
    .X(_05142_));
 sky130_fd_sc_hd__buf_1 _09657_ (.A(_05142_),
    .X(_05143_));
 sky130_fd_sc_hd__a22o_1 _09658_ (.A1(\r1.regblock[30][8] ),
    .A2(_05131_),
    .B1(_05143_),
    .B2(_05135_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_1 _09659_ (.A(_05141_),
    .X(_01987_));
 sky130_fd_sc_hd__buf_1 _09660_ (.A(_05130_),
    .X(_05144_));
 sky130_fd_sc_hd__buf_1 _09661_ (.A(_04563_),
    .X(_05145_));
 sky130_fd_sc_hd__buf_1 _09662_ (.A(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__buf_1 _09663_ (.A(_05134_),
    .X(_05147_));
 sky130_fd_sc_hd__a22o_1 _09664_ (.A1(\r1.regblock[30][7] ),
    .A2(_05144_),
    .B1(_05146_),
    .B2(_05147_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_1 _09665_ (.A(_05141_),
    .X(_01986_));
 sky130_fd_sc_hd__buf_1 _09666_ (.A(_04567_),
    .X(_05148_));
 sky130_fd_sc_hd__buf_1 _09667_ (.A(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__a22o_1 _09668_ (.A1(\r1.regblock[30][6] ),
    .A2(_05144_),
    .B1(_05149_),
    .B2(_05147_),
    .X(_03011_));
 sky130_fd_sc_hd__buf_1 _09669_ (.A(_05140_),
    .X(_05150_));
 sky130_fd_sc_hd__clkbuf_1 _09670_ (.A(_05150_),
    .X(_01985_));
 sky130_fd_sc_hd__buf_1 _09671_ (.A(_04571_),
    .X(_05151_));
 sky130_fd_sc_hd__buf_1 _09672_ (.A(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__a22o_1 _09673_ (.A1(\r1.regblock[30][5] ),
    .A2(_05144_),
    .B1(_05152_),
    .B2(_05147_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_1 _09674_ (.A(_05150_),
    .X(_01984_));
 sky130_fd_sc_hd__buf_1 _09675_ (.A(_05130_),
    .X(_05153_));
 sky130_fd_sc_hd__buf_1 _09676_ (.A(_04575_),
    .X(_05154_));
 sky130_fd_sc_hd__buf_1 _09677_ (.A(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__buf_1 _09678_ (.A(_05134_),
    .X(_05156_));
 sky130_fd_sc_hd__a22o_1 _09679_ (.A1(\r1.regblock[30][4] ),
    .A2(_05153_),
    .B1(_05155_),
    .B2(_05156_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_1 _09680_ (.A(_05150_),
    .X(_01983_));
 sky130_fd_sc_hd__buf_1 _09681_ (.A(_04579_),
    .X(_05157_));
 sky130_fd_sc_hd__buf_1 _09682_ (.A(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__a22o_1 _09683_ (.A1(\r1.regblock[30][3] ),
    .A2(_05153_),
    .B1(_05158_),
    .B2(_05156_),
    .X(_03008_));
 sky130_fd_sc_hd__buf_1 _09684_ (.A(_05140_),
    .X(_05159_));
 sky130_fd_sc_hd__clkbuf_1 _09685_ (.A(_05159_),
    .X(_01982_));
 sky130_fd_sc_hd__buf_1 _09686_ (.A(_04583_),
    .X(_05160_));
 sky130_fd_sc_hd__buf_1 _09687_ (.A(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__a22o_1 _09688_ (.A1(\r1.regblock[30][2] ),
    .A2(_05153_),
    .B1(_05161_),
    .B2(_05156_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_1 _09689_ (.A(_05159_),
    .X(_01981_));
 sky130_fd_sc_hd__buf_1 _09690_ (.A(_04586_),
    .X(_05162_));
 sky130_fd_sc_hd__buf_1 _09691_ (.A(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__a22o_1 _09692_ (.A1(\r1.regblock[30][1] ),
    .A2(_05056_),
    .B1(_05163_),
    .B2(_05061_),
    .X(_03006_));
 sky130_fd_sc_hd__clkbuf_1 _09693_ (.A(_05159_),
    .X(_01980_));
 sky130_fd_sc_hd__buf_1 _09694_ (.A(_04589_),
    .X(_05164_));
 sky130_fd_sc_hd__buf_1 _09695_ (.A(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__a22o_1 _09696_ (.A1(\r1.regblock[30][0] ),
    .A2(_05056_),
    .B1(_05165_),
    .B2(_05061_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_4 _09697_ (.A(_05139_),
    .X(_05166_));
 sky130_fd_sc_hd__buf_1 _09698_ (.A(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__clkbuf_1 _09699_ (.A(_05167_),
    .X(_01979_));
 sky130_fd_sc_hd__or2_2 _09700_ (.A(_04217_),
    .B(_05053_),
    .X(_05168_));
 sky130_fd_sc_hd__buf_1 _09701_ (.A(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__buf_1 _09702_ (.A(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__inv_2 _09703_ (.A(_05168_),
    .Y(_05171_));
 sky130_fd_sc_hd__buf_1 _09704_ (.A(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__buf_1 _09705_ (.A(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__a22o_1 _09706_ (.A1(\r1.regblock[2][31] ),
    .A2(_05170_),
    .B1(_05059_),
    .B2(_05173_),
    .X(_03004_));
 sky130_fd_sc_hd__clkbuf_1 _09707_ (.A(_05167_),
    .X(_01978_));
 sky130_fd_sc_hd__a22o_1 _09708_ (.A1(\r1.regblock[2][30] ),
    .A2(_05170_),
    .B1(_05064_),
    .B2(_05173_),
    .X(_03003_));
 sky130_fd_sc_hd__clkbuf_1 _09709_ (.A(_05167_),
    .X(_01977_));
 sky130_fd_sc_hd__a22o_1 _09710_ (.A1(\r1.regblock[2][29] ),
    .A2(_05170_),
    .B1(_05067_),
    .B2(_05173_),
    .X(_03002_));
 sky130_fd_sc_hd__buf_1 _09711_ (.A(_05166_),
    .X(_05174_));
 sky130_fd_sc_hd__clkbuf_1 _09712_ (.A(_05174_),
    .X(_01976_));
 sky130_fd_sc_hd__clkbuf_4 _09713_ (.A(_05168_),
    .X(_05175_));
 sky130_fd_sc_hd__clkbuf_2 _09714_ (.A(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__buf_1 _09715_ (.A(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__clkbuf_4 _09716_ (.A(_05171_),
    .X(_05178_));
 sky130_fd_sc_hd__clkbuf_2 _09717_ (.A(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__buf_1 _09718_ (.A(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__a22o_1 _09719_ (.A1(\r1.regblock[2][28] ),
    .A2(_05177_),
    .B1(_05072_),
    .B2(_05180_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_1 _09720_ (.A(_05174_),
    .X(_01975_));
 sky130_fd_sc_hd__a22o_1 _09721_ (.A1(\r1.regblock[2][27] ),
    .A2(_05177_),
    .B1(_05077_),
    .B2(_05180_),
    .X(_03000_));
 sky130_fd_sc_hd__clkbuf_1 _09722_ (.A(_05174_),
    .X(_01974_));
 sky130_fd_sc_hd__a22o_1 _09723_ (.A1(\r1.regblock[2][26] ),
    .A2(_05177_),
    .B1(_05081_),
    .B2(_05180_),
    .X(_02999_));
 sky130_fd_sc_hd__buf_1 _09724_ (.A(_05166_),
    .X(_05181_));
 sky130_fd_sc_hd__clkbuf_1 _09725_ (.A(_05181_),
    .X(_01973_));
 sky130_fd_sc_hd__buf_1 _09726_ (.A(_05176_),
    .X(_05182_));
 sky130_fd_sc_hd__buf_1 _09727_ (.A(_05179_),
    .X(_05183_));
 sky130_fd_sc_hd__a22o_1 _09728_ (.A1(\r1.regblock[2][25] ),
    .A2(_05182_),
    .B1(_05084_),
    .B2(_05183_),
    .X(_02998_));
 sky130_fd_sc_hd__clkbuf_1 _09729_ (.A(_05181_),
    .X(_01972_));
 sky130_fd_sc_hd__a22o_1 _09730_ (.A1(\r1.regblock[2][24] ),
    .A2(_05182_),
    .B1(_05087_),
    .B2(_05183_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_1 _09731_ (.A(_05181_),
    .X(_01971_));
 sky130_fd_sc_hd__a22o_1 _09732_ (.A1(\r1.regblock[2][23] ),
    .A2(_05182_),
    .B1(_05090_),
    .B2(_05183_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_4 _09733_ (.A(_05139_),
    .X(_05184_));
 sky130_fd_sc_hd__buf_1 _09734_ (.A(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__clkbuf_1 _09735_ (.A(_05185_),
    .X(_01970_));
 sky130_fd_sc_hd__buf_1 _09736_ (.A(_05176_),
    .X(_05186_));
 sky130_fd_sc_hd__buf_1 _09737_ (.A(_05179_),
    .X(_05187_));
 sky130_fd_sc_hd__a22o_1 _09738_ (.A1(\r1.regblock[2][22] ),
    .A2(_05186_),
    .B1(_05093_),
    .B2(_05187_),
    .X(_02995_));
 sky130_fd_sc_hd__clkbuf_1 _09739_ (.A(_05185_),
    .X(_01969_));
 sky130_fd_sc_hd__a22o_1 _09740_ (.A1(\r1.regblock[2][21] ),
    .A2(_05186_),
    .B1(_05096_),
    .B2(_05187_),
    .X(_02994_));
 sky130_fd_sc_hd__clkbuf_1 _09741_ (.A(_05185_),
    .X(_01968_));
 sky130_fd_sc_hd__a22o_1 _09742_ (.A1(\r1.regblock[2][20] ),
    .A2(_05186_),
    .B1(_05099_),
    .B2(_05187_),
    .X(_02993_));
 sky130_fd_sc_hd__clkbuf_1 _09743_ (.A(_05184_),
    .X(_05188_));
 sky130_fd_sc_hd__clkbuf_1 _09744_ (.A(_05188_),
    .X(_01967_));
 sky130_fd_sc_hd__clkbuf_2 _09745_ (.A(_05175_),
    .X(_05189_));
 sky130_fd_sc_hd__buf_1 _09746_ (.A(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__clkbuf_2 _09747_ (.A(_05178_),
    .X(_05191_));
 sky130_fd_sc_hd__buf_1 _09748_ (.A(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__a22o_1 _09749_ (.A1(\r1.regblock[2][19] ),
    .A2(_05190_),
    .B1(_05103_),
    .B2(_05192_),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _09750_ (.A(_05188_),
    .X(_01966_));
 sky130_fd_sc_hd__a22o_1 _09751_ (.A1(\r1.regblock[2][18] ),
    .A2(_05190_),
    .B1(_05107_),
    .B2(_05192_),
    .X(_02991_));
 sky130_fd_sc_hd__clkbuf_1 _09752_ (.A(_05188_),
    .X(_01965_));
 sky130_fd_sc_hd__a22o_1 _09753_ (.A1(\r1.regblock[2][17] ),
    .A2(_05190_),
    .B1(_05111_),
    .B2(_05192_),
    .X(_02990_));
 sky130_fd_sc_hd__buf_1 _09754_ (.A(_05184_),
    .X(_05193_));
 sky130_fd_sc_hd__clkbuf_1 _09755_ (.A(_05193_),
    .X(_01964_));
 sky130_fd_sc_hd__buf_1 _09756_ (.A(_05189_),
    .X(_05194_));
 sky130_fd_sc_hd__buf_1 _09757_ (.A(_05191_),
    .X(_05195_));
 sky130_fd_sc_hd__a22o_1 _09758_ (.A1(\r1.regblock[2][16] ),
    .A2(_05194_),
    .B1(_05114_),
    .B2(_05195_),
    .X(_02989_));
 sky130_fd_sc_hd__clkbuf_1 _09759_ (.A(_05193_),
    .X(_01963_));
 sky130_fd_sc_hd__a22o_1 _09760_ (.A1(\r1.regblock[2][15] ),
    .A2(_05194_),
    .B1(_05117_),
    .B2(_05195_),
    .X(_02988_));
 sky130_fd_sc_hd__clkbuf_1 _09761_ (.A(_05193_),
    .X(_01962_));
 sky130_fd_sc_hd__a22o_1 _09762_ (.A1(\r1.regblock[2][14] ),
    .A2(_05194_),
    .B1(_05120_),
    .B2(_05195_),
    .X(_02987_));
 sky130_fd_sc_hd__buf_1 _09763_ (.A(_05138_),
    .X(_05196_));
 sky130_fd_sc_hd__clkbuf_4 _09764_ (.A(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__buf_1 _09765_ (.A(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__clkbuf_1 _09766_ (.A(_05198_),
    .X(_01961_));
 sky130_fd_sc_hd__buf_1 _09767_ (.A(_05189_),
    .X(_05199_));
 sky130_fd_sc_hd__buf_1 _09768_ (.A(_05191_),
    .X(_05200_));
 sky130_fd_sc_hd__a22o_1 _09769_ (.A1(\r1.regblock[2][13] ),
    .A2(_05199_),
    .B1(_05123_),
    .B2(_05200_),
    .X(_02986_));
 sky130_fd_sc_hd__clkbuf_1 _09770_ (.A(_05198_),
    .X(_01960_));
 sky130_fd_sc_hd__a22o_1 _09771_ (.A1(\r1.regblock[2][12] ),
    .A2(_05199_),
    .B1(_05126_),
    .B2(_05200_),
    .X(_02985_));
 sky130_fd_sc_hd__clkbuf_1 _09772_ (.A(_05198_),
    .X(_01959_));
 sky130_fd_sc_hd__a22o_1 _09773_ (.A1(\r1.regblock[2][11] ),
    .A2(_05199_),
    .B1(_05129_),
    .B2(_05200_),
    .X(_02984_));
 sky130_fd_sc_hd__buf_1 _09774_ (.A(_05197_),
    .X(_05201_));
 sky130_fd_sc_hd__clkbuf_1 _09775_ (.A(_05201_),
    .X(_01958_));
 sky130_fd_sc_hd__buf_1 _09776_ (.A(_05175_),
    .X(_05202_));
 sky130_fd_sc_hd__buf_1 _09777_ (.A(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__buf_1 _09778_ (.A(_05178_),
    .X(_05204_));
 sky130_fd_sc_hd__buf_1 _09779_ (.A(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__a22o_1 _09780_ (.A1(\r1.regblock[2][10] ),
    .A2(_05203_),
    .B1(_05133_),
    .B2(_05205_),
    .X(_02983_));
 sky130_fd_sc_hd__clkbuf_1 _09781_ (.A(_05201_),
    .X(_01957_));
 sky130_fd_sc_hd__a22o_1 _09782_ (.A1(\r1.regblock[2][9] ),
    .A2(_05203_),
    .B1(_05137_),
    .B2(_05205_),
    .X(_02982_));
 sky130_fd_sc_hd__clkbuf_1 _09783_ (.A(_05201_),
    .X(_01956_));
 sky130_fd_sc_hd__a22o_1 _09784_ (.A1(\r1.regblock[2][8] ),
    .A2(_05203_),
    .B1(_05143_),
    .B2(_05205_),
    .X(_02981_));
 sky130_fd_sc_hd__buf_1 _09785_ (.A(_05197_),
    .X(_05206_));
 sky130_fd_sc_hd__clkbuf_1 _09786_ (.A(_05206_),
    .X(_01955_));
 sky130_fd_sc_hd__buf_1 _09787_ (.A(_05202_),
    .X(_05207_));
 sky130_fd_sc_hd__buf_1 _09788_ (.A(_05204_),
    .X(_05208_));
 sky130_fd_sc_hd__a22o_1 _09789_ (.A1(\r1.regblock[2][7] ),
    .A2(_05207_),
    .B1(_05146_),
    .B2(_05208_),
    .X(_02980_));
 sky130_fd_sc_hd__clkbuf_1 _09790_ (.A(_05206_),
    .X(_01954_));
 sky130_fd_sc_hd__a22o_1 _09791_ (.A1(\r1.regblock[2][6] ),
    .A2(_05207_),
    .B1(_05149_),
    .B2(_05208_),
    .X(_02979_));
 sky130_fd_sc_hd__clkbuf_1 _09792_ (.A(_05206_),
    .X(_01953_));
 sky130_fd_sc_hd__a22o_1 _09793_ (.A1(\r1.regblock[2][5] ),
    .A2(_05207_),
    .B1(_05152_),
    .B2(_05208_),
    .X(_02978_));
 sky130_fd_sc_hd__buf_2 _09794_ (.A(_05196_),
    .X(_05209_));
 sky130_fd_sc_hd__buf_1 _09795_ (.A(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__clkbuf_1 _09796_ (.A(_05210_),
    .X(_01952_));
 sky130_fd_sc_hd__buf_1 _09797_ (.A(_05202_),
    .X(_05211_));
 sky130_fd_sc_hd__buf_1 _09798_ (.A(_05204_),
    .X(_05212_));
 sky130_fd_sc_hd__a22o_1 _09799_ (.A1(\r1.regblock[2][4] ),
    .A2(_05211_),
    .B1(_05155_),
    .B2(_05212_),
    .X(_02977_));
 sky130_fd_sc_hd__clkbuf_1 _09800_ (.A(_05210_),
    .X(_01951_));
 sky130_fd_sc_hd__a22o_1 _09801_ (.A1(\r1.regblock[2][3] ),
    .A2(_05211_),
    .B1(_05158_),
    .B2(_05212_),
    .X(_02976_));
 sky130_fd_sc_hd__clkbuf_1 _09802_ (.A(_05210_),
    .X(_01950_));
 sky130_fd_sc_hd__a22o_1 _09803_ (.A1(\r1.regblock[2][2] ),
    .A2(_05211_),
    .B1(_05161_),
    .B2(_05212_),
    .X(_02975_));
 sky130_fd_sc_hd__buf_1 _09804_ (.A(_05209_),
    .X(_05213_));
 sky130_fd_sc_hd__clkbuf_1 _09805_ (.A(_05213_),
    .X(_01949_));
 sky130_fd_sc_hd__a22o_1 _09806_ (.A1(\r1.regblock[2][1] ),
    .A2(_05169_),
    .B1(_05163_),
    .B2(_05172_),
    .X(_02974_));
 sky130_fd_sc_hd__clkbuf_1 _09807_ (.A(_05213_),
    .X(_01948_));
 sky130_fd_sc_hd__a22o_1 _09808_ (.A1(\r1.regblock[2][0] ),
    .A2(_05169_),
    .B1(_05165_),
    .B2(_05172_),
    .X(_02973_));
 sky130_fd_sc_hd__clkbuf_1 _09809_ (.A(_05213_),
    .X(_01947_));
 sky130_fd_sc_hd__or2_2 _09810_ (.A(_04776_),
    .B(_04954_),
    .X(_05214_));
 sky130_fd_sc_hd__buf_1 _09811_ (.A(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__buf_1 _09812_ (.A(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__inv_2 _09813_ (.A(_05214_),
    .Y(_05217_));
 sky130_fd_sc_hd__buf_1 _09814_ (.A(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__buf_1 _09815_ (.A(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__a22o_1 _09816_ (.A1(\r1.regblock[28][31] ),
    .A2(_05216_),
    .B1(_05059_),
    .B2(_05219_),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_2 _09817_ (.A(_05209_),
    .X(_05220_));
 sky130_fd_sc_hd__clkbuf_1 _09818_ (.A(_05220_),
    .X(_01946_));
 sky130_fd_sc_hd__a22o_1 _09819_ (.A1(\r1.regblock[28][30] ),
    .A2(_05216_),
    .B1(_05064_),
    .B2(_05219_),
    .X(_02971_));
 sky130_fd_sc_hd__clkbuf_1 _09820_ (.A(_05220_),
    .X(_01945_));
 sky130_fd_sc_hd__a22o_1 _09821_ (.A1(\r1.regblock[28][29] ),
    .A2(_05216_),
    .B1(_05067_),
    .B2(_05219_),
    .X(_02970_));
 sky130_fd_sc_hd__clkbuf_1 _09822_ (.A(_05220_),
    .X(_01944_));
 sky130_fd_sc_hd__clkbuf_4 _09823_ (.A(_05214_),
    .X(_05221_));
 sky130_fd_sc_hd__buf_2 _09824_ (.A(_05221_),
    .X(_05222_));
 sky130_fd_sc_hd__buf_1 _09825_ (.A(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__buf_2 _09826_ (.A(_05217_),
    .X(_05224_));
 sky130_fd_sc_hd__buf_2 _09827_ (.A(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__buf_1 _09828_ (.A(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__a22o_1 _09829_ (.A1(\r1.regblock[28][28] ),
    .A2(_05223_),
    .B1(_05072_),
    .B2(_05226_),
    .X(_02969_));
 sky130_fd_sc_hd__clkbuf_2 _09830_ (.A(_05196_),
    .X(_05227_));
 sky130_fd_sc_hd__clkbuf_2 _09831_ (.A(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__clkbuf_1 _09832_ (.A(_05228_),
    .X(_01943_));
 sky130_fd_sc_hd__a22o_1 _09833_ (.A1(\r1.regblock[28][27] ),
    .A2(_05223_),
    .B1(_05077_),
    .B2(_05226_),
    .X(_02968_));
 sky130_fd_sc_hd__clkbuf_1 _09834_ (.A(_05228_),
    .X(_01942_));
 sky130_fd_sc_hd__a22o_1 _09835_ (.A1(\r1.regblock[28][26] ),
    .A2(_05223_),
    .B1(_05081_),
    .B2(_05226_),
    .X(_02967_));
 sky130_fd_sc_hd__clkbuf_1 _09836_ (.A(_05228_),
    .X(_01941_));
 sky130_fd_sc_hd__buf_1 _09837_ (.A(_05222_),
    .X(_05229_));
 sky130_fd_sc_hd__buf_1 _09838_ (.A(_05225_),
    .X(_05230_));
 sky130_fd_sc_hd__a22o_1 _09839_ (.A1(\r1.regblock[28][25] ),
    .A2(_05229_),
    .B1(_05084_),
    .B2(_05230_),
    .X(_02966_));
 sky130_fd_sc_hd__buf_1 _09840_ (.A(_05227_),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_1 _09841_ (.A(_05231_),
    .X(_01940_));
 sky130_fd_sc_hd__a22o_1 _09842_ (.A1(\r1.regblock[28][24] ),
    .A2(_05229_),
    .B1(_05087_),
    .B2(_05230_),
    .X(_02965_));
 sky130_fd_sc_hd__clkbuf_1 _09843_ (.A(_05231_),
    .X(_01939_));
 sky130_fd_sc_hd__a22o_1 _09844_ (.A1(\r1.regblock[28][23] ),
    .A2(_05229_),
    .B1(_05090_),
    .B2(_05230_),
    .X(_02964_));
 sky130_fd_sc_hd__clkbuf_1 _09845_ (.A(_05231_),
    .X(_01938_));
 sky130_fd_sc_hd__buf_1 _09846_ (.A(_05222_),
    .X(_05232_));
 sky130_fd_sc_hd__buf_1 _09847_ (.A(_05225_),
    .X(_05233_));
 sky130_fd_sc_hd__a22o_1 _09848_ (.A1(\r1.regblock[28][22] ),
    .A2(_05232_),
    .B1(_05093_),
    .B2(_05233_),
    .X(_02963_));
 sky130_fd_sc_hd__buf_1 _09849_ (.A(_05227_),
    .X(_05234_));
 sky130_fd_sc_hd__clkbuf_1 _09850_ (.A(_05234_),
    .X(_01937_));
 sky130_fd_sc_hd__a22o_1 _09851_ (.A1(\r1.regblock[28][21] ),
    .A2(_05232_),
    .B1(_05096_),
    .B2(_05233_),
    .X(_02962_));
 sky130_fd_sc_hd__clkbuf_1 _09852_ (.A(_05234_),
    .X(_01936_));
 sky130_fd_sc_hd__a22o_1 _09853_ (.A1(\r1.regblock[28][20] ),
    .A2(_05232_),
    .B1(_05099_),
    .B2(_05233_),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_2 _09854_ (.A(_05234_),
    .X(_01935_));
 sky130_fd_sc_hd__clkbuf_2 _09855_ (.A(_05221_),
    .X(_05235_));
 sky130_fd_sc_hd__buf_1 _09856_ (.A(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__buf_2 _09857_ (.A(_05224_),
    .X(_05237_));
 sky130_fd_sc_hd__buf_1 _09858_ (.A(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__a22o_1 _09859_ (.A1(\r1.regblock[28][19] ),
    .A2(_05236_),
    .B1(_05103_),
    .B2(_05238_),
    .X(_02960_));
 sky130_fd_sc_hd__buf_2 _09860_ (.A(_05138_),
    .X(_05239_));
 sky130_fd_sc_hd__clkbuf_4 _09861_ (.A(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__buf_1 _09862_ (.A(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__clkbuf_1 _09863_ (.A(_05241_),
    .X(_01934_));
 sky130_fd_sc_hd__a22o_1 _09864_ (.A1(\r1.regblock[28][18] ),
    .A2(_05236_),
    .B1(_05107_),
    .B2(_05238_),
    .X(_02959_));
 sky130_fd_sc_hd__clkbuf_1 _09865_ (.A(_05241_),
    .X(_01933_));
 sky130_fd_sc_hd__a22o_1 _09866_ (.A1(\r1.regblock[28][17] ),
    .A2(_05236_),
    .B1(_05111_),
    .B2(_05238_),
    .X(_02958_));
 sky130_fd_sc_hd__clkbuf_1 _09867_ (.A(_05241_),
    .X(_01932_));
 sky130_fd_sc_hd__buf_1 _09868_ (.A(_05235_),
    .X(_05242_));
 sky130_fd_sc_hd__buf_1 _09869_ (.A(_05237_),
    .X(_05243_));
 sky130_fd_sc_hd__a22o_1 _09870_ (.A1(\r1.regblock[28][16] ),
    .A2(_05242_),
    .B1(_05114_),
    .B2(_05243_),
    .X(_02957_));
 sky130_fd_sc_hd__buf_1 _09871_ (.A(_05240_),
    .X(_05244_));
 sky130_fd_sc_hd__clkbuf_1 _09872_ (.A(_05244_),
    .X(_01931_));
 sky130_fd_sc_hd__a22o_1 _09873_ (.A1(\r1.regblock[28][15] ),
    .A2(_05242_),
    .B1(_05117_),
    .B2(_05243_),
    .X(_02956_));
 sky130_fd_sc_hd__clkbuf_1 _09874_ (.A(_05244_),
    .X(_01930_));
 sky130_fd_sc_hd__a22o_1 _09875_ (.A1(\r1.regblock[28][14] ),
    .A2(_05242_),
    .B1(_05120_),
    .B2(_05243_),
    .X(_02955_));
 sky130_fd_sc_hd__clkbuf_1 _09876_ (.A(_05244_),
    .X(_01929_));
 sky130_fd_sc_hd__buf_1 _09877_ (.A(_05235_),
    .X(_05245_));
 sky130_fd_sc_hd__buf_1 _09878_ (.A(_05237_),
    .X(_05246_));
 sky130_fd_sc_hd__a22o_1 _09879_ (.A1(\r1.regblock[28][13] ),
    .A2(_05245_),
    .B1(_05123_),
    .B2(_05246_),
    .X(_02954_));
 sky130_fd_sc_hd__buf_2 _09880_ (.A(_05240_),
    .X(_05247_));
 sky130_fd_sc_hd__clkbuf_1 _09881_ (.A(_05247_),
    .X(_01928_));
 sky130_fd_sc_hd__a22o_1 _09882_ (.A1(\r1.regblock[28][12] ),
    .A2(_05245_),
    .B1(_05126_),
    .B2(_05246_),
    .X(_02953_));
 sky130_fd_sc_hd__clkbuf_1 _09883_ (.A(_05247_),
    .X(_01927_));
 sky130_fd_sc_hd__a22o_1 _09884_ (.A1(\r1.regblock[28][11] ),
    .A2(_05245_),
    .B1(_05129_),
    .B2(_05246_),
    .X(_02952_));
 sky130_fd_sc_hd__clkbuf_1 _09885_ (.A(_05247_),
    .X(_01926_));
 sky130_fd_sc_hd__clkbuf_2 _09886_ (.A(_05221_),
    .X(_05248_));
 sky130_fd_sc_hd__buf_1 _09887_ (.A(_05248_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_2 _09888_ (.A(_05224_),
    .X(_05250_));
 sky130_fd_sc_hd__buf_1 _09889_ (.A(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__a22o_1 _09890_ (.A1(\r1.regblock[28][10] ),
    .A2(_05249_),
    .B1(_05133_),
    .B2(_05251_),
    .X(_02951_));
 sky130_fd_sc_hd__buf_1 _09891_ (.A(_05239_),
    .X(_05252_));
 sky130_fd_sc_hd__buf_1 _09892_ (.A(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__clkbuf_1 _09893_ (.A(_05253_),
    .X(_01925_));
 sky130_fd_sc_hd__a22o_1 _09894_ (.A1(\r1.regblock[28][9] ),
    .A2(_05249_),
    .B1(_05137_),
    .B2(_05251_),
    .X(_02950_));
 sky130_fd_sc_hd__clkbuf_1 _09895_ (.A(_05253_),
    .X(_01924_));
 sky130_fd_sc_hd__a22o_1 _09896_ (.A1(\r1.regblock[28][8] ),
    .A2(_05249_),
    .B1(_05143_),
    .B2(_05251_),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_1 _09897_ (.A(_05253_),
    .X(_01923_));
 sky130_fd_sc_hd__buf_1 _09898_ (.A(_05248_),
    .X(_05254_));
 sky130_fd_sc_hd__buf_1 _09899_ (.A(_05250_),
    .X(_05255_));
 sky130_fd_sc_hd__a22o_1 _09900_ (.A1(\r1.regblock[28][7] ),
    .A2(_05254_),
    .B1(_05146_),
    .B2(_05255_),
    .X(_02948_));
 sky130_fd_sc_hd__buf_1 _09901_ (.A(_05252_),
    .X(_05256_));
 sky130_fd_sc_hd__clkbuf_1 _09902_ (.A(_05256_),
    .X(_01922_));
 sky130_fd_sc_hd__a22o_1 _09903_ (.A1(\r1.regblock[28][6] ),
    .A2(_05254_),
    .B1(_05149_),
    .B2(_05255_),
    .X(_02947_));
 sky130_fd_sc_hd__clkbuf_1 _09904_ (.A(_05256_),
    .X(_01921_));
 sky130_fd_sc_hd__a22o_1 _09905_ (.A1(\r1.regblock[28][5] ),
    .A2(_05254_),
    .B1(_05152_),
    .B2(_05255_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_1 _09906_ (.A(_05256_),
    .X(_01920_));
 sky130_fd_sc_hd__buf_1 _09907_ (.A(_05248_),
    .X(_05257_));
 sky130_fd_sc_hd__buf_1 _09908_ (.A(_05250_),
    .X(_05258_));
 sky130_fd_sc_hd__a22o_1 _09909_ (.A1(\r1.regblock[28][4] ),
    .A2(_05257_),
    .B1(_05155_),
    .B2(_05258_),
    .X(_02945_));
 sky130_fd_sc_hd__buf_1 _09910_ (.A(_05252_),
    .X(_05259_));
 sky130_fd_sc_hd__clkbuf_1 _09911_ (.A(_05259_),
    .X(_01919_));
 sky130_fd_sc_hd__a22o_1 _09912_ (.A1(\r1.regblock[28][3] ),
    .A2(_05257_),
    .B1(_05158_),
    .B2(_05258_),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_1 _09913_ (.A(_05259_),
    .X(_01918_));
 sky130_fd_sc_hd__a22o_1 _09914_ (.A1(\r1.regblock[28][2] ),
    .A2(_05257_),
    .B1(_05161_),
    .B2(_05258_),
    .X(_02943_));
 sky130_fd_sc_hd__buf_1 _09915_ (.A(_05259_),
    .X(_01917_));
 sky130_fd_sc_hd__a22o_1 _09916_ (.A1(\r1.regblock[28][1] ),
    .A2(_05215_),
    .B1(_05163_),
    .B2(_05218_),
    .X(_02942_));
 sky130_fd_sc_hd__buf_1 _09917_ (.A(_05239_),
    .X(_05260_));
 sky130_fd_sc_hd__buf_1 _09918_ (.A(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__clkbuf_1 _09919_ (.A(_05261_),
    .X(_01916_));
 sky130_fd_sc_hd__a22o_1 _09920_ (.A1(\r1.regblock[28][0] ),
    .A2(_05215_),
    .B1(_05165_),
    .B2(_05218_),
    .X(_02941_));
 sky130_fd_sc_hd__clkbuf_1 _09921_ (.A(_05261_),
    .X(_01915_));
 sky130_fd_sc_hd__buf_1 _09922_ (.A(_04223_),
    .X(_05262_));
 sky130_fd_sc_hd__or3_1 _09923_ (.A(_04341_),
    .B(_04389_),
    .C(\r1.waddr[2] ),
    .X(_05263_));
 sky130_fd_sc_hd__clkbuf_1 _09924_ (.A(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__or2_2 _09925_ (.A(_05262_),
    .B(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__buf_1 _09926_ (.A(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__buf_1 _09927_ (.A(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__buf_1 _09928_ (.A(_05058_),
    .X(_05268_));
 sky130_fd_sc_hd__inv_2 _09929_ (.A(_05265_),
    .Y(_05269_));
 sky130_fd_sc_hd__buf_1 _09930_ (.A(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__buf_1 _09931_ (.A(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__a22o_1 _09932_ (.A1(\r1.regblock[27][31] ),
    .A2(_05267_),
    .B1(_05268_),
    .B2(_05271_),
    .X(_02940_));
 sky130_fd_sc_hd__clkbuf_1 _09933_ (.A(_05261_),
    .X(_01914_));
 sky130_fd_sc_hd__buf_1 _09934_ (.A(_05063_),
    .X(_05272_));
 sky130_fd_sc_hd__a22o_1 _09935_ (.A1(\r1.regblock[27][30] ),
    .A2(_05267_),
    .B1(_05272_),
    .B2(_05271_),
    .X(_02939_));
 sky130_fd_sc_hd__buf_1 _09936_ (.A(_05260_),
    .X(_05273_));
 sky130_fd_sc_hd__clkbuf_1 _09937_ (.A(_05273_),
    .X(_01913_));
 sky130_fd_sc_hd__buf_1 _09938_ (.A(_05066_),
    .X(_05274_));
 sky130_fd_sc_hd__a22o_1 _09939_ (.A1(\r1.regblock[27][29] ),
    .A2(_05267_),
    .B1(_05274_),
    .B2(_05271_),
    .X(_02938_));
 sky130_fd_sc_hd__clkbuf_1 _09940_ (.A(_05273_),
    .X(_01912_));
 sky130_fd_sc_hd__clkbuf_2 _09941_ (.A(_05265_),
    .X(_05275_));
 sky130_fd_sc_hd__buf_2 _09942_ (.A(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__buf_1 _09943_ (.A(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__buf_1 _09944_ (.A(_05071_),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_2 _09945_ (.A(_05269_),
    .X(_05279_));
 sky130_fd_sc_hd__buf_2 _09946_ (.A(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__buf_1 _09947_ (.A(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__a22o_1 _09948_ (.A1(\r1.regblock[27][28] ),
    .A2(_05277_),
    .B1(_05278_),
    .B2(_05281_),
    .X(_02937_));
 sky130_fd_sc_hd__clkbuf_1 _09949_ (.A(_05273_),
    .X(_01911_));
 sky130_fd_sc_hd__buf_1 _09950_ (.A(_05076_),
    .X(_05282_));
 sky130_fd_sc_hd__a22o_1 _09951_ (.A1(\r1.regblock[27][27] ),
    .A2(_05277_),
    .B1(_05282_),
    .B2(_05281_),
    .X(_02936_));
 sky130_fd_sc_hd__buf_1 _09952_ (.A(_05260_),
    .X(_05283_));
 sky130_fd_sc_hd__clkbuf_1 _09953_ (.A(_05283_),
    .X(_01910_));
 sky130_fd_sc_hd__buf_1 _09954_ (.A(_05080_),
    .X(_05284_));
 sky130_fd_sc_hd__a22o_1 _09955_ (.A1(\r1.regblock[27][26] ),
    .A2(_05277_),
    .B1(_05284_),
    .B2(_05281_),
    .X(_02935_));
 sky130_fd_sc_hd__clkbuf_1 _09956_ (.A(_05283_),
    .X(_01909_));
 sky130_fd_sc_hd__buf_1 _09957_ (.A(_05276_),
    .X(_05285_));
 sky130_fd_sc_hd__buf_1 _09958_ (.A(_05083_),
    .X(_05286_));
 sky130_fd_sc_hd__buf_1 _09959_ (.A(_05280_),
    .X(_05287_));
 sky130_fd_sc_hd__a22o_1 _09960_ (.A1(\r1.regblock[27][25] ),
    .A2(_05285_),
    .B1(_05286_),
    .B2(_05287_),
    .X(_02934_));
 sky130_fd_sc_hd__clkbuf_1 _09961_ (.A(_05283_),
    .X(_01908_));
 sky130_fd_sc_hd__buf_1 _09962_ (.A(_05086_),
    .X(_05288_));
 sky130_fd_sc_hd__a22o_1 _09963_ (.A1(\r1.regblock[27][24] ),
    .A2(_05285_),
    .B1(_05288_),
    .B2(_05287_),
    .X(_02933_));
 sky130_fd_sc_hd__buf_1 _09964_ (.A(_04969_),
    .X(_05289_));
 sky130_fd_sc_hd__clkbuf_2 _09965_ (.A(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__buf_2 _09966_ (.A(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__buf_1 _09967_ (.A(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__buf_1 _09968_ (.A(_05292_),
    .X(_01907_));
 sky130_fd_sc_hd__buf_1 _09969_ (.A(_05089_),
    .X(_05293_));
 sky130_fd_sc_hd__a22o_1 _09970_ (.A1(\r1.regblock[27][23] ),
    .A2(_05285_),
    .B1(_05293_),
    .B2(_05287_),
    .X(_02932_));
 sky130_fd_sc_hd__clkbuf_1 _09971_ (.A(_05292_),
    .X(_01906_));
 sky130_fd_sc_hd__buf_1 _09972_ (.A(_05276_),
    .X(_05294_));
 sky130_fd_sc_hd__buf_1 _09973_ (.A(_05092_),
    .X(_05295_));
 sky130_fd_sc_hd__buf_1 _09974_ (.A(_05280_),
    .X(_05296_));
 sky130_fd_sc_hd__a22o_1 _09975_ (.A1(\r1.regblock[27][22] ),
    .A2(_05294_),
    .B1(_05295_),
    .B2(_05296_),
    .X(_02931_));
 sky130_fd_sc_hd__clkbuf_1 _09976_ (.A(_05292_),
    .X(_01905_));
 sky130_fd_sc_hd__buf_1 _09977_ (.A(_05095_),
    .X(_05297_));
 sky130_fd_sc_hd__a22o_1 _09978_ (.A1(\r1.regblock[27][21] ),
    .A2(_05294_),
    .B1(_05297_),
    .B2(_05296_),
    .X(_02930_));
 sky130_fd_sc_hd__buf_1 _09979_ (.A(_05291_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_2 _09980_ (.A(_05298_),
    .X(_01904_));
 sky130_fd_sc_hd__buf_1 _09981_ (.A(_05098_),
    .X(_05299_));
 sky130_fd_sc_hd__a22o_1 _09982_ (.A1(\r1.regblock[27][20] ),
    .A2(_05294_),
    .B1(_05299_),
    .B2(_05296_),
    .X(_02929_));
 sky130_fd_sc_hd__clkbuf_1 _09983_ (.A(_05298_),
    .X(_01903_));
 sky130_fd_sc_hd__buf_2 _09984_ (.A(_05275_),
    .X(_05300_));
 sky130_fd_sc_hd__buf_1 _09985_ (.A(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__buf_1 _09986_ (.A(_05102_),
    .X(_05302_));
 sky130_fd_sc_hd__buf_2 _09987_ (.A(_05279_),
    .X(_05303_));
 sky130_fd_sc_hd__buf_1 _09988_ (.A(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__a22o_1 _09989_ (.A1(\r1.regblock[27][19] ),
    .A2(_05301_),
    .B1(_05302_),
    .B2(_05304_),
    .X(_02928_));
 sky130_fd_sc_hd__clkbuf_1 _09990_ (.A(_05298_),
    .X(_01902_));
 sky130_fd_sc_hd__buf_1 _09991_ (.A(_05106_),
    .X(_05305_));
 sky130_fd_sc_hd__a22o_1 _09992_ (.A1(\r1.regblock[27][18] ),
    .A2(_05301_),
    .B1(_05305_),
    .B2(_05304_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_2 _09993_ (.A(_05291_),
    .X(_05306_));
 sky130_fd_sc_hd__clkbuf_1 _09994_ (.A(_05306_),
    .X(_01901_));
 sky130_fd_sc_hd__buf_1 _09995_ (.A(_05110_),
    .X(_05307_));
 sky130_fd_sc_hd__a22o_1 _09996_ (.A1(\r1.regblock[27][17] ),
    .A2(_05301_),
    .B1(_05307_),
    .B2(_05304_),
    .X(_02926_));
 sky130_fd_sc_hd__clkbuf_1 _09997_ (.A(_05306_),
    .X(_01900_));
 sky130_fd_sc_hd__buf_1 _09998_ (.A(_05300_),
    .X(_05308_));
 sky130_fd_sc_hd__buf_1 _09999_ (.A(_05113_),
    .X(_05309_));
 sky130_fd_sc_hd__buf_1 _10000_ (.A(_05303_),
    .X(_05310_));
 sky130_fd_sc_hd__a22o_1 _10001_ (.A1(\r1.regblock[27][16] ),
    .A2(_05308_),
    .B1(_05309_),
    .B2(_05310_),
    .X(_02925_));
 sky130_fd_sc_hd__clkbuf_1 _10002_ (.A(_05306_),
    .X(_01899_));
 sky130_fd_sc_hd__buf_1 _10003_ (.A(_05116_),
    .X(_05311_));
 sky130_fd_sc_hd__a22o_1 _10004_ (.A1(\r1.regblock[27][15] ),
    .A2(_05308_),
    .B1(_05311_),
    .B2(_05310_),
    .X(_02924_));
 sky130_fd_sc_hd__buf_2 _10005_ (.A(_05290_),
    .X(_05312_));
 sky130_fd_sc_hd__buf_1 _10006_ (.A(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__clkbuf_1 _10007_ (.A(_05313_),
    .X(_01898_));
 sky130_fd_sc_hd__buf_1 _10008_ (.A(_05119_),
    .X(_05314_));
 sky130_fd_sc_hd__a22o_1 _10009_ (.A1(\r1.regblock[27][14] ),
    .A2(_05308_),
    .B1(_05314_),
    .B2(_05310_),
    .X(_02923_));
 sky130_fd_sc_hd__clkbuf_1 _10010_ (.A(_05313_),
    .X(_01897_));
 sky130_fd_sc_hd__buf_1 _10011_ (.A(_05300_),
    .X(_05315_));
 sky130_fd_sc_hd__buf_1 _10012_ (.A(_05122_),
    .X(_05316_));
 sky130_fd_sc_hd__buf_1 _10013_ (.A(_05303_),
    .X(_05317_));
 sky130_fd_sc_hd__a22o_1 _10014_ (.A1(\r1.regblock[27][13] ),
    .A2(_05315_),
    .B1(_05316_),
    .B2(_05317_),
    .X(_02922_));
 sky130_fd_sc_hd__clkbuf_1 _10015_ (.A(_05313_),
    .X(_01896_));
 sky130_fd_sc_hd__buf_1 _10016_ (.A(_05125_),
    .X(_05318_));
 sky130_fd_sc_hd__a22o_1 _10017_ (.A1(\r1.regblock[27][12] ),
    .A2(_05315_),
    .B1(_05318_),
    .B2(_05317_),
    .X(_02921_));
 sky130_fd_sc_hd__clkbuf_2 _10018_ (.A(_05312_),
    .X(_05319_));
 sky130_fd_sc_hd__clkbuf_1 _10019_ (.A(_05319_),
    .X(_01895_));
 sky130_fd_sc_hd__buf_1 _10020_ (.A(_05128_),
    .X(_05320_));
 sky130_fd_sc_hd__a22o_1 _10021_ (.A1(\r1.regblock[27][11] ),
    .A2(_05315_),
    .B1(_05320_),
    .B2(_05317_),
    .X(_02920_));
 sky130_fd_sc_hd__clkbuf_1 _10022_ (.A(_05319_),
    .X(_01894_));
 sky130_fd_sc_hd__clkbuf_2 _10023_ (.A(_05275_),
    .X(_05321_));
 sky130_fd_sc_hd__buf_1 _10024_ (.A(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__buf_1 _10025_ (.A(_05132_),
    .X(_05323_));
 sky130_fd_sc_hd__clkbuf_2 _10026_ (.A(_05279_),
    .X(_05324_));
 sky130_fd_sc_hd__buf_1 _10027_ (.A(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__a22o_1 _10028_ (.A1(\r1.regblock[27][10] ),
    .A2(_05322_),
    .B1(_05323_),
    .B2(_05325_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_1 _10029_ (.A(_05319_),
    .X(_01893_));
 sky130_fd_sc_hd__buf_1 _10030_ (.A(_05136_),
    .X(_05326_));
 sky130_fd_sc_hd__a22o_1 _10031_ (.A1(\r1.regblock[27][9] ),
    .A2(_05322_),
    .B1(_05326_),
    .B2(_05325_),
    .X(_02918_));
 sky130_fd_sc_hd__buf_1 _10032_ (.A(_05312_),
    .X(_05327_));
 sky130_fd_sc_hd__clkbuf_1 _10033_ (.A(_05327_),
    .X(_01892_));
 sky130_fd_sc_hd__buf_1 _10034_ (.A(_05142_),
    .X(_05328_));
 sky130_fd_sc_hd__a22o_1 _10035_ (.A1(\r1.regblock[27][8] ),
    .A2(_05322_),
    .B1(_05328_),
    .B2(_05325_),
    .X(_02917_));
 sky130_fd_sc_hd__clkbuf_1 _10036_ (.A(_05327_),
    .X(_01891_));
 sky130_fd_sc_hd__buf_1 _10037_ (.A(_05321_),
    .X(_05329_));
 sky130_fd_sc_hd__buf_1 _10038_ (.A(_05145_),
    .X(_05330_));
 sky130_fd_sc_hd__buf_1 _10039_ (.A(_05324_),
    .X(_05331_));
 sky130_fd_sc_hd__a22o_1 _10040_ (.A1(\r1.regblock[27][7] ),
    .A2(_05329_),
    .B1(_05330_),
    .B2(_05331_),
    .X(_02916_));
 sky130_fd_sc_hd__clkbuf_1 _10041_ (.A(_05327_),
    .X(_01890_));
 sky130_fd_sc_hd__buf_1 _10042_ (.A(_05148_),
    .X(_05332_));
 sky130_fd_sc_hd__a22o_1 _10043_ (.A1(\r1.regblock[27][6] ),
    .A2(_05329_),
    .B1(_05332_),
    .B2(_05331_),
    .X(_02915_));
 sky130_fd_sc_hd__clkbuf_2 _10044_ (.A(_05290_),
    .X(_05333_));
 sky130_fd_sc_hd__buf_1 _10045_ (.A(_05333_),
    .X(_05334_));
 sky130_fd_sc_hd__buf_1 _10046_ (.A(_05334_),
    .X(_01889_));
 sky130_fd_sc_hd__buf_1 _10047_ (.A(_05151_),
    .X(_05335_));
 sky130_fd_sc_hd__a22o_1 _10048_ (.A1(\r1.regblock[27][5] ),
    .A2(_05329_),
    .B1(_05335_),
    .B2(_05331_),
    .X(_02914_));
 sky130_fd_sc_hd__clkbuf_1 _10049_ (.A(_05334_),
    .X(_01888_));
 sky130_fd_sc_hd__buf_1 _10050_ (.A(_05321_),
    .X(_05336_));
 sky130_fd_sc_hd__buf_1 _10051_ (.A(_05154_),
    .X(_05337_));
 sky130_fd_sc_hd__buf_1 _10052_ (.A(_05324_),
    .X(_05338_));
 sky130_fd_sc_hd__a22o_1 _10053_ (.A1(\r1.regblock[27][4] ),
    .A2(_05336_),
    .B1(_05337_),
    .B2(_05338_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_1 _10054_ (.A(_05334_),
    .X(_01887_));
 sky130_fd_sc_hd__buf_1 _10055_ (.A(_05157_),
    .X(_05339_));
 sky130_fd_sc_hd__a22o_1 _10056_ (.A1(\r1.regblock[27][3] ),
    .A2(_05336_),
    .B1(_05339_),
    .B2(_05338_),
    .X(_02912_));
 sky130_fd_sc_hd__buf_1 _10057_ (.A(_05333_),
    .X(_05340_));
 sky130_fd_sc_hd__clkbuf_1 _10058_ (.A(_05340_),
    .X(_01886_));
 sky130_fd_sc_hd__buf_1 _10059_ (.A(_05160_),
    .X(_05341_));
 sky130_fd_sc_hd__a22o_1 _10060_ (.A1(\r1.regblock[27][2] ),
    .A2(_05336_),
    .B1(_05341_),
    .B2(_05338_),
    .X(_02911_));
 sky130_fd_sc_hd__clkbuf_1 _10061_ (.A(_05340_),
    .X(_01885_));
 sky130_fd_sc_hd__buf_1 _10062_ (.A(_05162_),
    .X(_05342_));
 sky130_fd_sc_hd__a22o_1 _10063_ (.A1(\r1.regblock[27][1] ),
    .A2(_05266_),
    .B1(_05342_),
    .B2(_05270_),
    .X(_02910_));
 sky130_fd_sc_hd__clkbuf_1 _10064_ (.A(_05340_),
    .X(_01884_));
 sky130_fd_sc_hd__buf_1 _10065_ (.A(_05164_),
    .X(_05343_));
 sky130_fd_sc_hd__a22o_1 _10066_ (.A1(\r1.regblock[27][0] ),
    .A2(_05266_),
    .B1(_05343_),
    .B2(_05270_),
    .X(_02909_));
 sky130_fd_sc_hd__buf_1 _10067_ (.A(_05333_),
    .X(_05344_));
 sky130_fd_sc_hd__clkbuf_1 _10068_ (.A(_05344_),
    .X(_01883_));
 sky130_fd_sc_hd__or2_2 _10069_ (.A(_05054_),
    .B(_05264_),
    .X(_05345_));
 sky130_fd_sc_hd__buf_1 _10070_ (.A(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__buf_1 _10071_ (.A(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__inv_2 _10072_ (.A(_05345_),
    .Y(_05348_));
 sky130_fd_sc_hd__buf_1 _10073_ (.A(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__buf_1 _10074_ (.A(_05349_),
    .X(_05350_));
 sky130_fd_sc_hd__a22o_1 _10075_ (.A1(\r1.regblock[26][31] ),
    .A2(_05347_),
    .B1(_05268_),
    .B2(_05350_),
    .X(_02908_));
 sky130_fd_sc_hd__clkbuf_1 _10076_ (.A(_05344_),
    .X(_01882_));
 sky130_fd_sc_hd__a22o_1 _10077_ (.A1(\r1.regblock[26][30] ),
    .A2(_05347_),
    .B1(_05272_),
    .B2(_05350_),
    .X(_02907_));
 sky130_fd_sc_hd__clkbuf_1 _10078_ (.A(_05344_),
    .X(_01881_));
 sky130_fd_sc_hd__a22o_1 _10079_ (.A1(\r1.regblock[26][29] ),
    .A2(_05347_),
    .B1(_05274_),
    .B2(_05350_),
    .X(_02906_));
 sky130_fd_sc_hd__buf_1 _10080_ (.A(_05289_),
    .X(_05351_));
 sky130_fd_sc_hd__buf_2 _10081_ (.A(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__buf_1 _10082_ (.A(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__clkbuf_1 _10083_ (.A(_05353_),
    .X(_01880_));
 sky130_fd_sc_hd__clkbuf_2 _10084_ (.A(_05345_),
    .X(_05354_));
 sky130_fd_sc_hd__buf_2 _10085_ (.A(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__buf_1 _10086_ (.A(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__clkbuf_2 _10087_ (.A(_05348_),
    .X(_05357_));
 sky130_fd_sc_hd__buf_2 _10088_ (.A(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__buf_1 _10089_ (.A(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__a22o_1 _10090_ (.A1(\r1.regblock[26][28] ),
    .A2(_05356_),
    .B1(_05278_),
    .B2(_05359_),
    .X(_02905_));
 sky130_fd_sc_hd__clkbuf_1 _10091_ (.A(_05353_),
    .X(_01879_));
 sky130_fd_sc_hd__a22o_1 _10092_ (.A1(\r1.regblock[26][27] ),
    .A2(_05356_),
    .B1(_05282_),
    .B2(_05359_),
    .X(_02904_));
 sky130_fd_sc_hd__clkbuf_1 _10093_ (.A(_05353_),
    .X(_01878_));
 sky130_fd_sc_hd__a22o_1 _10094_ (.A1(\r1.regblock[26][26] ),
    .A2(_05356_),
    .B1(_05284_),
    .B2(_05359_),
    .X(_02903_));
 sky130_fd_sc_hd__buf_1 _10095_ (.A(_05352_),
    .X(_05360_));
 sky130_fd_sc_hd__clkbuf_1 _10096_ (.A(_05360_),
    .X(_01877_));
 sky130_fd_sc_hd__buf_1 _10097_ (.A(_05355_),
    .X(_05361_));
 sky130_fd_sc_hd__buf_1 _10098_ (.A(_05358_),
    .X(_05362_));
 sky130_fd_sc_hd__a22o_1 _10099_ (.A1(\r1.regblock[26][25] ),
    .A2(_05361_),
    .B1(_05286_),
    .B2(_05362_),
    .X(_02902_));
 sky130_fd_sc_hd__clkbuf_1 _10100_ (.A(_05360_),
    .X(_01876_));
 sky130_fd_sc_hd__a22o_1 _10101_ (.A1(\r1.regblock[26][24] ),
    .A2(_05361_),
    .B1(_05288_),
    .B2(_05362_),
    .X(_02901_));
 sky130_fd_sc_hd__clkbuf_1 _10102_ (.A(_05360_),
    .X(_01875_));
 sky130_fd_sc_hd__a22o_1 _10103_ (.A1(\r1.regblock[26][23] ),
    .A2(_05361_),
    .B1(_05293_),
    .B2(_05362_),
    .X(_02900_));
 sky130_fd_sc_hd__buf_1 _10104_ (.A(_05352_),
    .X(_05363_));
 sky130_fd_sc_hd__clkbuf_1 _10105_ (.A(_05363_),
    .X(_01874_));
 sky130_fd_sc_hd__buf_1 _10106_ (.A(_05355_),
    .X(_05364_));
 sky130_fd_sc_hd__buf_1 _10107_ (.A(_05358_),
    .X(_05365_));
 sky130_fd_sc_hd__a22o_1 _10108_ (.A1(\r1.regblock[26][22] ),
    .A2(_05364_),
    .B1(_05295_),
    .B2(_05365_),
    .X(_02899_));
 sky130_fd_sc_hd__clkbuf_1 _10109_ (.A(_05363_),
    .X(_01873_));
 sky130_fd_sc_hd__a22o_1 _10110_ (.A1(\r1.regblock[26][21] ),
    .A2(_05364_),
    .B1(_05297_),
    .B2(_05365_),
    .X(_02898_));
 sky130_fd_sc_hd__clkbuf_1 _10111_ (.A(_05363_),
    .X(_01872_));
 sky130_fd_sc_hd__a22o_1 _10112_ (.A1(\r1.regblock[26][20] ),
    .A2(_05364_),
    .B1(_05299_),
    .B2(_05365_),
    .X(_02897_));
 sky130_fd_sc_hd__clkbuf_4 _10113_ (.A(_05351_),
    .X(_05366_));
 sky130_fd_sc_hd__buf_1 _10114_ (.A(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__clkbuf_1 _10115_ (.A(_05367_),
    .X(_01871_));
 sky130_fd_sc_hd__buf_2 _10116_ (.A(_05354_),
    .X(_05368_));
 sky130_fd_sc_hd__buf_1 _10117_ (.A(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__buf_2 _10118_ (.A(_05357_),
    .X(_05370_));
 sky130_fd_sc_hd__buf_1 _10119_ (.A(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__a22o_1 _10120_ (.A1(\r1.regblock[26][19] ),
    .A2(_05369_),
    .B1(_05302_),
    .B2(_05371_),
    .X(_02896_));
 sky130_fd_sc_hd__clkbuf_1 _10121_ (.A(_05367_),
    .X(_01870_));
 sky130_fd_sc_hd__a22o_1 _10122_ (.A1(\r1.regblock[26][18] ),
    .A2(_05369_),
    .B1(_05305_),
    .B2(_05371_),
    .X(_02895_));
 sky130_fd_sc_hd__clkbuf_1 _10123_ (.A(_05367_),
    .X(_01869_));
 sky130_fd_sc_hd__a22o_1 _10124_ (.A1(\r1.regblock[26][17] ),
    .A2(_05369_),
    .B1(_05307_),
    .B2(_05371_),
    .X(_02894_));
 sky130_fd_sc_hd__buf_1 _10125_ (.A(_05366_),
    .X(_05372_));
 sky130_fd_sc_hd__clkbuf_1 _10126_ (.A(_05372_),
    .X(_01868_));
 sky130_fd_sc_hd__buf_1 _10127_ (.A(_05368_),
    .X(_05373_));
 sky130_fd_sc_hd__buf_1 _10128_ (.A(_05370_),
    .X(_05374_));
 sky130_fd_sc_hd__a22o_1 _10129_ (.A1(\r1.regblock[26][16] ),
    .A2(_05373_),
    .B1(_05309_),
    .B2(_05374_),
    .X(_02893_));
 sky130_fd_sc_hd__clkbuf_1 _10130_ (.A(_05372_),
    .X(_01867_));
 sky130_fd_sc_hd__a22o_1 _10131_ (.A1(\r1.regblock[26][15] ),
    .A2(_05373_),
    .B1(_05311_),
    .B2(_05374_),
    .X(_02892_));
 sky130_fd_sc_hd__clkbuf_1 _10132_ (.A(_05372_),
    .X(_01866_));
 sky130_fd_sc_hd__a22o_1 _10133_ (.A1(\r1.regblock[26][14] ),
    .A2(_05373_),
    .B1(_05314_),
    .B2(_05374_),
    .X(_02891_));
 sky130_fd_sc_hd__buf_1 _10134_ (.A(_05366_),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_1 _10135_ (.A(_05375_),
    .X(_01865_));
 sky130_fd_sc_hd__buf_1 _10136_ (.A(_05368_),
    .X(_05376_));
 sky130_fd_sc_hd__buf_1 _10137_ (.A(_05370_),
    .X(_05377_));
 sky130_fd_sc_hd__a22o_1 _10138_ (.A1(\r1.regblock[26][13] ),
    .A2(_05376_),
    .B1(_05316_),
    .B2(_05377_),
    .X(_02890_));
 sky130_fd_sc_hd__clkbuf_1 _10139_ (.A(_05375_),
    .X(_01864_));
 sky130_fd_sc_hd__a22o_1 _10140_ (.A1(\r1.regblock[26][12] ),
    .A2(_05376_),
    .B1(_05318_),
    .B2(_05377_),
    .X(_02889_));
 sky130_fd_sc_hd__clkbuf_1 _10141_ (.A(_05375_),
    .X(_01863_));
 sky130_fd_sc_hd__a22o_1 _10142_ (.A1(\r1.regblock[26][11] ),
    .A2(_05376_),
    .B1(_05320_),
    .B2(_05377_),
    .X(_02888_));
 sky130_fd_sc_hd__clkbuf_2 _10143_ (.A(_05351_),
    .X(_05378_));
 sky130_fd_sc_hd__buf_1 _10144_ (.A(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__clkbuf_1 _10145_ (.A(_05379_),
    .X(_01862_));
 sky130_fd_sc_hd__clkbuf_2 _10146_ (.A(_05354_),
    .X(_05380_));
 sky130_fd_sc_hd__buf_1 _10147_ (.A(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__clkbuf_2 _10148_ (.A(_05357_),
    .X(_05382_));
 sky130_fd_sc_hd__buf_1 _10149_ (.A(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__a22o_1 _10150_ (.A1(\r1.regblock[26][10] ),
    .A2(_05381_),
    .B1(_05323_),
    .B2(_05383_),
    .X(_02887_));
 sky130_fd_sc_hd__clkbuf_1 _10151_ (.A(_05379_),
    .X(_01861_));
 sky130_fd_sc_hd__a22o_1 _10152_ (.A1(\r1.regblock[26][9] ),
    .A2(_05381_),
    .B1(_05326_),
    .B2(_05383_),
    .X(_02886_));
 sky130_fd_sc_hd__clkbuf_1 _10153_ (.A(_05379_),
    .X(_01860_));
 sky130_fd_sc_hd__a22o_1 _10154_ (.A1(\r1.regblock[26][8] ),
    .A2(_05381_),
    .B1(_05328_),
    .B2(_05383_),
    .X(_02885_));
 sky130_fd_sc_hd__buf_1 _10155_ (.A(_05378_),
    .X(_05384_));
 sky130_fd_sc_hd__clkbuf_1 _10156_ (.A(_05384_),
    .X(_01859_));
 sky130_fd_sc_hd__buf_1 _10157_ (.A(_05380_),
    .X(_05385_));
 sky130_fd_sc_hd__buf_1 _10158_ (.A(_05382_),
    .X(_05386_));
 sky130_fd_sc_hd__a22o_1 _10159_ (.A1(\r1.regblock[26][7] ),
    .A2(_05385_),
    .B1(_05330_),
    .B2(_05386_),
    .X(_02884_));
 sky130_fd_sc_hd__clkbuf_1 _10160_ (.A(_05384_),
    .X(_01858_));
 sky130_fd_sc_hd__a22o_1 _10161_ (.A1(\r1.regblock[26][6] ),
    .A2(_05385_),
    .B1(_05332_),
    .B2(_05386_),
    .X(_02883_));
 sky130_fd_sc_hd__clkbuf_1 _10162_ (.A(_05384_),
    .X(_01857_));
 sky130_fd_sc_hd__a22o_1 _10163_ (.A1(\r1.regblock[26][5] ),
    .A2(_05385_),
    .B1(_05335_),
    .B2(_05386_),
    .X(_02882_));
 sky130_fd_sc_hd__buf_1 _10164_ (.A(_05378_),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _10165_ (.A(_05387_),
    .X(_01856_));
 sky130_fd_sc_hd__buf_1 _10166_ (.A(_05380_),
    .X(_05388_));
 sky130_fd_sc_hd__buf_1 _10167_ (.A(_05382_),
    .X(_05389_));
 sky130_fd_sc_hd__a22o_1 _10168_ (.A1(\r1.regblock[26][4] ),
    .A2(_05388_),
    .B1(_05337_),
    .B2(_05389_),
    .X(_02881_));
 sky130_fd_sc_hd__clkbuf_1 _10169_ (.A(_05387_),
    .X(_01855_));
 sky130_fd_sc_hd__a22o_1 _10170_ (.A1(\r1.regblock[26][3] ),
    .A2(_05388_),
    .B1(_05339_),
    .B2(_05389_),
    .X(_02880_));
 sky130_fd_sc_hd__clkbuf_1 _10171_ (.A(_05387_),
    .X(_01854_));
 sky130_fd_sc_hd__a22o_1 _10172_ (.A1(\r1.regblock[26][2] ),
    .A2(_05388_),
    .B1(_05341_),
    .B2(_05389_),
    .X(_02879_));
 sky130_fd_sc_hd__buf_1 _10173_ (.A(_05289_),
    .X(_05390_));
 sky130_fd_sc_hd__buf_2 _10174_ (.A(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__buf_1 _10175_ (.A(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__clkbuf_1 _10176_ (.A(_05392_),
    .X(_01853_));
 sky130_fd_sc_hd__a22o_1 _10177_ (.A1(\r1.regblock[26][1] ),
    .A2(_05346_),
    .B1(_05342_),
    .B2(_05349_),
    .X(_02878_));
 sky130_fd_sc_hd__clkbuf_1 _10178_ (.A(_05392_),
    .X(_01852_));
 sky130_fd_sc_hd__a22o_1 _10179_ (.A1(\r1.regblock[26][0] ),
    .A2(_05346_),
    .B1(_05343_),
    .B2(_05349_),
    .X(_02877_));
 sky130_fd_sc_hd__clkbuf_1 _10180_ (.A(_05392_),
    .X(_01851_));
 sky130_fd_sc_hd__or2_2 _10181_ (.A(_04396_),
    .B(_05264_),
    .X(_05393_));
 sky130_fd_sc_hd__buf_1 _10182_ (.A(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__buf_1 _10183_ (.A(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__inv_2 _10184_ (.A(_05393_),
    .Y(_05396_));
 sky130_fd_sc_hd__buf_1 _10185_ (.A(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__buf_1 _10186_ (.A(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__a22o_1 _10187_ (.A1(\r1.regblock[25][31] ),
    .A2(_05395_),
    .B1(_05268_),
    .B2(_05398_),
    .X(_02876_));
 sky130_fd_sc_hd__buf_1 _10188_ (.A(_05391_),
    .X(_05399_));
 sky130_fd_sc_hd__clkbuf_1 _10189_ (.A(_05399_),
    .X(_01850_));
 sky130_fd_sc_hd__a22o_1 _10190_ (.A1(\r1.regblock[25][30] ),
    .A2(_05395_),
    .B1(_05272_),
    .B2(_05398_),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_1 _10191_ (.A(_05399_),
    .X(_01849_));
 sky130_fd_sc_hd__a22o_1 _10192_ (.A1(\r1.regblock[25][29] ),
    .A2(_05395_),
    .B1(_05274_),
    .B2(_05398_),
    .X(_02874_));
 sky130_fd_sc_hd__clkbuf_1 _10193_ (.A(_05399_),
    .X(_01848_));
 sky130_fd_sc_hd__clkbuf_2 _10194_ (.A(_05393_),
    .X(_05400_));
 sky130_fd_sc_hd__buf_2 _10195_ (.A(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__buf_1 _10196_ (.A(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_2 _10197_ (.A(_05396_),
    .X(_05403_));
 sky130_fd_sc_hd__buf_2 _10198_ (.A(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__buf_1 _10199_ (.A(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__a22o_1 _10200_ (.A1(\r1.regblock[25][28] ),
    .A2(_05402_),
    .B1(_05278_),
    .B2(_05405_),
    .X(_02873_));
 sky130_fd_sc_hd__buf_1 _10201_ (.A(_05391_),
    .X(_05406_));
 sky130_fd_sc_hd__clkbuf_1 _10202_ (.A(_05406_),
    .X(_01847_));
 sky130_fd_sc_hd__a22o_1 _10203_ (.A1(\r1.regblock[25][27] ),
    .A2(_05402_),
    .B1(_05282_),
    .B2(_05405_),
    .X(_02872_));
 sky130_fd_sc_hd__clkbuf_1 _10204_ (.A(_05406_),
    .X(_01846_));
 sky130_fd_sc_hd__a22o_1 _10205_ (.A1(\r1.regblock[25][26] ),
    .A2(_05402_),
    .B1(_05284_),
    .B2(_05405_),
    .X(_02871_));
 sky130_fd_sc_hd__clkbuf_1 _10206_ (.A(_05406_),
    .X(_01845_));
 sky130_fd_sc_hd__buf_1 _10207_ (.A(_05401_),
    .X(_05407_));
 sky130_fd_sc_hd__buf_1 _10208_ (.A(_05404_),
    .X(_05408_));
 sky130_fd_sc_hd__a22o_1 _10209_ (.A1(\r1.regblock[25][25] ),
    .A2(_05407_),
    .B1(_05286_),
    .B2(_05408_),
    .X(_02870_));
 sky130_fd_sc_hd__buf_1 _10210_ (.A(_05390_),
    .X(_05409_));
 sky130_fd_sc_hd__clkbuf_2 _10211_ (.A(_05409_),
    .X(_05410_));
 sky130_fd_sc_hd__clkbuf_1 _10212_ (.A(_05410_),
    .X(_01844_));
 sky130_fd_sc_hd__a22o_1 _10213_ (.A1(\r1.regblock[25][24] ),
    .A2(_05407_),
    .B1(_05288_),
    .B2(_05408_),
    .X(_02869_));
 sky130_fd_sc_hd__clkbuf_1 _10214_ (.A(_05410_),
    .X(_01843_));
 sky130_fd_sc_hd__a22o_1 _10215_ (.A1(\r1.regblock[25][23] ),
    .A2(_05407_),
    .B1(_05293_),
    .B2(_05408_),
    .X(_02868_));
 sky130_fd_sc_hd__clkbuf_1 _10216_ (.A(_05410_),
    .X(_01842_));
 sky130_fd_sc_hd__buf_1 _10217_ (.A(_05401_),
    .X(_05411_));
 sky130_fd_sc_hd__buf_1 _10218_ (.A(_05404_),
    .X(_05412_));
 sky130_fd_sc_hd__a22o_1 _10219_ (.A1(\r1.regblock[25][22] ),
    .A2(_05411_),
    .B1(_05295_),
    .B2(_05412_),
    .X(_02867_));
 sky130_fd_sc_hd__buf_2 _10220_ (.A(_05409_),
    .X(_05413_));
 sky130_fd_sc_hd__clkbuf_1 _10221_ (.A(_05413_),
    .X(_01841_));
 sky130_fd_sc_hd__a22o_1 _10222_ (.A1(\r1.regblock[25][21] ),
    .A2(_05411_),
    .B1(_05297_),
    .B2(_05412_),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_1 _10223_ (.A(_05413_),
    .X(_01840_));
 sky130_fd_sc_hd__a22o_1 _10224_ (.A1(\r1.regblock[25][20] ),
    .A2(_05411_),
    .B1(_05299_),
    .B2(_05412_),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_1 _10225_ (.A(_05413_),
    .X(_01839_));
 sky130_fd_sc_hd__buf_2 _10226_ (.A(_05400_),
    .X(_05414_));
 sky130_fd_sc_hd__buf_1 _10227_ (.A(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__buf_2 _10228_ (.A(_05403_),
    .X(_05416_));
 sky130_fd_sc_hd__buf_1 _10229_ (.A(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__a22o_1 _10230_ (.A1(\r1.regblock[25][19] ),
    .A2(_05415_),
    .B1(_05302_),
    .B2(_05417_),
    .X(_02864_));
 sky130_fd_sc_hd__buf_2 _10231_ (.A(_05409_),
    .X(_05418_));
 sky130_fd_sc_hd__clkbuf_1 _10232_ (.A(_05418_),
    .X(_01838_));
 sky130_fd_sc_hd__a22o_1 _10233_ (.A1(\r1.regblock[25][18] ),
    .A2(_05415_),
    .B1(_05305_),
    .B2(_05417_),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _10234_ (.A(_05418_),
    .X(_01837_));
 sky130_fd_sc_hd__a22o_1 _10235_ (.A1(\r1.regblock[25][17] ),
    .A2(_05415_),
    .B1(_05307_),
    .B2(_05417_),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_1 _10236_ (.A(_05418_),
    .X(_01836_));
 sky130_fd_sc_hd__buf_1 _10237_ (.A(_05414_),
    .X(_05419_));
 sky130_fd_sc_hd__buf_1 _10238_ (.A(_05416_),
    .X(_05420_));
 sky130_fd_sc_hd__a22o_1 _10239_ (.A1(\r1.regblock[25][16] ),
    .A2(_05419_),
    .B1(_05309_),
    .B2(_05420_),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_4 _10240_ (.A(_05390_),
    .X(_05421_));
 sky130_fd_sc_hd__buf_1 _10241_ (.A(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__clkbuf_1 _10242_ (.A(_05422_),
    .X(_01835_));
 sky130_fd_sc_hd__a22o_1 _10243_ (.A1(\r1.regblock[25][15] ),
    .A2(_05419_),
    .B1(_05311_),
    .B2(_05420_),
    .X(_02860_));
 sky130_fd_sc_hd__clkbuf_1 _10244_ (.A(_05422_),
    .X(_01834_));
 sky130_fd_sc_hd__a22o_1 _10245_ (.A1(\r1.regblock[25][14] ),
    .A2(_05419_),
    .B1(_05314_),
    .B2(_05420_),
    .X(_02859_));
 sky130_fd_sc_hd__clkbuf_1 _10246_ (.A(_05422_),
    .X(_01833_));
 sky130_fd_sc_hd__buf_1 _10247_ (.A(_05414_),
    .X(_05423_));
 sky130_fd_sc_hd__buf_1 _10248_ (.A(_05416_),
    .X(_05424_));
 sky130_fd_sc_hd__a22o_1 _10249_ (.A1(\r1.regblock[25][13] ),
    .A2(_05423_),
    .B1(_05316_),
    .B2(_05424_),
    .X(_02858_));
 sky130_fd_sc_hd__clkbuf_2 _10250_ (.A(_05421_),
    .X(_05425_));
 sky130_fd_sc_hd__clkbuf_1 _10251_ (.A(_05425_),
    .X(_01832_));
 sky130_fd_sc_hd__a22o_1 _10252_ (.A1(\r1.regblock[25][12] ),
    .A2(_05423_),
    .B1(_05318_),
    .B2(_05424_),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _10253_ (.A(_05425_),
    .X(_01831_));
 sky130_fd_sc_hd__a22o_1 _10254_ (.A1(\r1.regblock[25][11] ),
    .A2(_05423_),
    .B1(_05320_),
    .B2(_05424_),
    .X(_02856_));
 sky130_fd_sc_hd__buf_1 _10255_ (.A(_05425_),
    .X(_01830_));
 sky130_fd_sc_hd__clkbuf_2 _10256_ (.A(_05400_),
    .X(_05426_));
 sky130_fd_sc_hd__buf_1 _10257_ (.A(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__clkbuf_2 _10258_ (.A(_05403_),
    .X(_05428_));
 sky130_fd_sc_hd__buf_1 _10259_ (.A(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__a22o_1 _10260_ (.A1(\r1.regblock[25][10] ),
    .A2(_05427_),
    .B1(_05323_),
    .B2(_05429_),
    .X(_02855_));
 sky130_fd_sc_hd__buf_1 _10261_ (.A(_05421_),
    .X(_05430_));
 sky130_fd_sc_hd__clkbuf_1 _10262_ (.A(_05430_),
    .X(_01829_));
 sky130_fd_sc_hd__a22o_1 _10263_ (.A1(\r1.regblock[25][9] ),
    .A2(_05427_),
    .B1(_05326_),
    .B2(_05429_),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _10264_ (.A(_05430_),
    .X(_01828_));
 sky130_fd_sc_hd__a22o_1 _10265_ (.A1(\r1.regblock[25][8] ),
    .A2(_05427_),
    .B1(_05328_),
    .B2(_05429_),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _10266_ (.A(_05430_),
    .X(_01827_));
 sky130_fd_sc_hd__buf_1 _10267_ (.A(_05426_),
    .X(_05431_));
 sky130_fd_sc_hd__buf_1 _10268_ (.A(_05428_),
    .X(_05432_));
 sky130_fd_sc_hd__a22o_1 _10269_ (.A1(\r1.regblock[25][7] ),
    .A2(_05431_),
    .B1(_05330_),
    .B2(_05432_),
    .X(_02852_));
 sky130_fd_sc_hd__buf_1 _10270_ (.A(_04429_),
    .X(_05433_));
 sky130_fd_sc_hd__buf_1 _10271_ (.A(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__buf_1 _10272_ (.A(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__buf_1 _10273_ (.A(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__clkbuf_2 _10274_ (.A(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__clkbuf_1 _10275_ (.A(_05437_),
    .X(_01826_));
 sky130_fd_sc_hd__a22o_1 _10276_ (.A1(\r1.regblock[25][6] ),
    .A2(_05431_),
    .B1(_05332_),
    .B2(_05432_),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _10277_ (.A(_05437_),
    .X(_01825_));
 sky130_fd_sc_hd__a22o_1 _10278_ (.A1(\r1.regblock[25][5] ),
    .A2(_05431_),
    .B1(_05335_),
    .B2(_05432_),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _10279_ (.A(_05437_),
    .X(_01824_));
 sky130_fd_sc_hd__buf_1 _10280_ (.A(_05426_),
    .X(_05438_));
 sky130_fd_sc_hd__buf_1 _10281_ (.A(_05428_),
    .X(_05439_));
 sky130_fd_sc_hd__a22o_1 _10282_ (.A1(\r1.regblock[25][4] ),
    .A2(_05438_),
    .B1(_05337_),
    .B2(_05439_),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_2 _10283_ (.A(_05436_),
    .X(_05440_));
 sky130_fd_sc_hd__clkbuf_1 _10284_ (.A(_05440_),
    .X(_01823_));
 sky130_fd_sc_hd__a22o_1 _10285_ (.A1(\r1.regblock[25][3] ),
    .A2(_05438_),
    .B1(_05339_),
    .B2(_05439_),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _10286_ (.A(_05440_),
    .X(_01822_));
 sky130_fd_sc_hd__a22o_1 _10287_ (.A1(\r1.regblock[25][2] ),
    .A2(_05438_),
    .B1(_05341_),
    .B2(_05439_),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _10288_ (.A(_05440_),
    .X(_01821_));
 sky130_fd_sc_hd__a22o_1 _10289_ (.A1(\r1.regblock[25][1] ),
    .A2(_05394_),
    .B1(_05342_),
    .B2(_05397_),
    .X(_02846_));
 sky130_fd_sc_hd__clkbuf_2 _10290_ (.A(_05436_),
    .X(_05441_));
 sky130_fd_sc_hd__clkbuf_1 _10291_ (.A(_05441_),
    .X(_01820_));
 sky130_fd_sc_hd__a22o_1 _10292_ (.A1(\r1.regblock[25][0] ),
    .A2(_05394_),
    .B1(_05343_),
    .B2(_05397_),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _10293_ (.A(_05441_),
    .X(_01819_));
 sky130_fd_sc_hd__or2_1 _10294_ (.A(_04776_),
    .B(_05263_),
    .X(_05442_));
 sky130_fd_sc_hd__buf_1 _10295_ (.A(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__buf_1 _10296_ (.A(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__buf_1 _10297_ (.A(_05058_),
    .X(_05445_));
 sky130_fd_sc_hd__inv_2 _10298_ (.A(_05442_),
    .Y(_05446_));
 sky130_fd_sc_hd__buf_1 _10299_ (.A(_05446_),
    .X(_05447_));
 sky130_fd_sc_hd__buf_1 _10300_ (.A(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__a22o_1 _10301_ (.A1(\r1.regblock[24][31] ),
    .A2(_05444_),
    .B1(_05445_),
    .B2(_05448_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _10302_ (.A(_05441_),
    .X(_01818_));
 sky130_fd_sc_hd__buf_1 _10303_ (.A(_05063_),
    .X(_05449_));
 sky130_fd_sc_hd__a22o_1 _10304_ (.A1(\r1.regblock[24][30] ),
    .A2(_05444_),
    .B1(_05449_),
    .B2(_05448_),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_2 _10305_ (.A(_05435_),
    .X(_05450_));
 sky130_fd_sc_hd__clkbuf_2 _10306_ (.A(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__clkbuf_1 _10307_ (.A(_05451_),
    .X(_01817_));
 sky130_fd_sc_hd__buf_1 _10308_ (.A(_05066_),
    .X(_05452_));
 sky130_fd_sc_hd__a22o_1 _10309_ (.A1(\r1.regblock[24][29] ),
    .A2(_05444_),
    .B1(_05452_),
    .B2(_05448_),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _10310_ (.A(_05451_),
    .X(_01816_));
 sky130_fd_sc_hd__buf_2 _10311_ (.A(_05442_),
    .X(_05453_));
 sky130_fd_sc_hd__buf_2 _10312_ (.A(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__buf_1 _10313_ (.A(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__clkbuf_2 _10314_ (.A(_05071_),
    .X(_05456_));
 sky130_fd_sc_hd__buf_2 _10315_ (.A(_05446_),
    .X(_05457_));
 sky130_fd_sc_hd__buf_2 _10316_ (.A(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__buf_1 _10317_ (.A(_05458_),
    .X(_05459_));
 sky130_fd_sc_hd__a22o_1 _10318_ (.A1(\r1.regblock[24][28] ),
    .A2(_05455_),
    .B1(_05456_),
    .B2(_05459_),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_1 _10319_ (.A(_05451_),
    .X(_01815_));
 sky130_fd_sc_hd__clkbuf_2 _10320_ (.A(_05076_),
    .X(_05460_));
 sky130_fd_sc_hd__a22o_1 _10321_ (.A1(\r1.regblock[24][27] ),
    .A2(_05455_),
    .B1(_05460_),
    .B2(_05459_),
    .X(_02840_));
 sky130_fd_sc_hd__buf_1 _10322_ (.A(_05450_),
    .X(_05461_));
 sky130_fd_sc_hd__clkbuf_1 _10323_ (.A(_05461_),
    .X(_01814_));
 sky130_fd_sc_hd__clkbuf_2 _10324_ (.A(_05080_),
    .X(_05462_));
 sky130_fd_sc_hd__a22o_1 _10325_ (.A1(\r1.regblock[24][26] ),
    .A2(_05455_),
    .B1(_05462_),
    .B2(_05459_),
    .X(_02839_));
 sky130_fd_sc_hd__clkbuf_1 _10326_ (.A(_05461_),
    .X(_01813_));
 sky130_fd_sc_hd__buf_1 _10327_ (.A(_05454_),
    .X(_05463_));
 sky130_fd_sc_hd__buf_1 _10328_ (.A(_05083_),
    .X(_05464_));
 sky130_fd_sc_hd__buf_1 _10329_ (.A(_05458_),
    .X(_05465_));
 sky130_fd_sc_hd__a22o_1 _10330_ (.A1(\r1.regblock[24][25] ),
    .A2(_05463_),
    .B1(_05464_),
    .B2(_05465_),
    .X(_02838_));
 sky130_fd_sc_hd__clkbuf_1 _10331_ (.A(_05461_),
    .X(_01812_));
 sky130_fd_sc_hd__buf_1 _10332_ (.A(_05086_),
    .X(_05466_));
 sky130_fd_sc_hd__a22o_1 _10333_ (.A1(\r1.regblock[24][24] ),
    .A2(_05463_),
    .B1(_05466_),
    .B2(_05465_),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_2 _10334_ (.A(_05450_),
    .X(_05467_));
 sky130_fd_sc_hd__clkbuf_1 _10335_ (.A(_05467_),
    .X(_01811_));
 sky130_fd_sc_hd__buf_1 _10336_ (.A(_05089_),
    .X(_05468_));
 sky130_fd_sc_hd__a22o_1 _10337_ (.A1(\r1.regblock[24][23] ),
    .A2(_05463_),
    .B1(_05468_),
    .B2(_05465_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _10338_ (.A(_05467_),
    .X(_01810_));
 sky130_fd_sc_hd__buf_1 _10339_ (.A(_05454_),
    .X(_05469_));
 sky130_fd_sc_hd__buf_1 _10340_ (.A(_05092_),
    .X(_05470_));
 sky130_fd_sc_hd__buf_1 _10341_ (.A(_05458_),
    .X(_05471_));
 sky130_fd_sc_hd__a22o_1 _10342_ (.A1(\r1.regblock[24][22] ),
    .A2(_05469_),
    .B1(_05470_),
    .B2(_05471_),
    .X(_02835_));
 sky130_fd_sc_hd__clkbuf_1 _10343_ (.A(_05467_),
    .X(_01809_));
 sky130_fd_sc_hd__buf_1 _10344_ (.A(_05095_),
    .X(_05472_));
 sky130_fd_sc_hd__a22o_1 _10345_ (.A1(\r1.regblock[24][21] ),
    .A2(_05469_),
    .B1(_05472_),
    .B2(_05471_),
    .X(_02834_));
 sky130_fd_sc_hd__buf_2 _10346_ (.A(_05435_),
    .X(_05473_));
 sky130_fd_sc_hd__buf_1 _10347_ (.A(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__clkbuf_2 _10348_ (.A(_05474_),
    .X(_01808_));
 sky130_fd_sc_hd__buf_1 _10349_ (.A(_05098_),
    .X(_05475_));
 sky130_fd_sc_hd__a22o_1 _10350_ (.A1(\r1.regblock[24][20] ),
    .A2(_05469_),
    .B1(_05475_),
    .B2(_05471_),
    .X(_02833_));
 sky130_fd_sc_hd__clkbuf_1 _10351_ (.A(_05474_),
    .X(_01807_));
 sky130_fd_sc_hd__buf_2 _10352_ (.A(_05453_),
    .X(_05476_));
 sky130_fd_sc_hd__buf_1 _10353_ (.A(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__clkbuf_2 _10354_ (.A(_05102_),
    .X(_05478_));
 sky130_fd_sc_hd__buf_2 _10355_ (.A(_05457_),
    .X(_05479_));
 sky130_fd_sc_hd__buf_1 _10356_ (.A(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__a22o_1 _10357_ (.A1(\r1.regblock[24][19] ),
    .A2(_05477_),
    .B1(_05478_),
    .B2(_05480_),
    .X(_02832_));
 sky130_fd_sc_hd__clkbuf_1 _10358_ (.A(_05474_),
    .X(_01806_));
 sky130_fd_sc_hd__clkbuf_2 _10359_ (.A(_05106_),
    .X(_05481_));
 sky130_fd_sc_hd__a22o_1 _10360_ (.A1(\r1.regblock[24][18] ),
    .A2(_05477_),
    .B1(_05481_),
    .B2(_05480_),
    .X(_02831_));
 sky130_fd_sc_hd__buf_1 _10361_ (.A(_05473_),
    .X(_05482_));
 sky130_fd_sc_hd__buf_1 _10362_ (.A(_05482_),
    .X(_01805_));
 sky130_fd_sc_hd__clkbuf_2 _10363_ (.A(_05110_),
    .X(_05483_));
 sky130_fd_sc_hd__a22o_1 _10364_ (.A1(\r1.regblock[24][17] ),
    .A2(_05477_),
    .B1(_05483_),
    .B2(_05480_),
    .X(_02830_));
 sky130_fd_sc_hd__clkbuf_1 _10365_ (.A(_05482_),
    .X(_01804_));
 sky130_fd_sc_hd__buf_1 _10366_ (.A(_05476_),
    .X(_05484_));
 sky130_fd_sc_hd__buf_1 _10367_ (.A(_05113_),
    .X(_05485_));
 sky130_fd_sc_hd__buf_1 _10368_ (.A(_05479_),
    .X(_05486_));
 sky130_fd_sc_hd__a22o_1 _10369_ (.A1(\r1.regblock[24][16] ),
    .A2(_05484_),
    .B1(_05485_),
    .B2(_05486_),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_1 _10370_ (.A(_05482_),
    .X(_01803_));
 sky130_fd_sc_hd__buf_1 _10371_ (.A(_05116_),
    .X(_05487_));
 sky130_fd_sc_hd__a22o_1 _10372_ (.A1(\r1.regblock[24][15] ),
    .A2(_05484_),
    .B1(_05487_),
    .B2(_05486_),
    .X(_02828_));
 sky130_fd_sc_hd__buf_1 _10373_ (.A(_05473_),
    .X(_05488_));
 sky130_fd_sc_hd__clkbuf_1 _10374_ (.A(_05488_),
    .X(_01802_));
 sky130_fd_sc_hd__buf_1 _10375_ (.A(_05119_),
    .X(_05489_));
 sky130_fd_sc_hd__a22o_1 _10376_ (.A1(\r1.regblock[24][14] ),
    .A2(_05484_),
    .B1(_05489_),
    .B2(_05486_),
    .X(_02827_));
 sky130_fd_sc_hd__clkbuf_1 _10377_ (.A(_05488_),
    .X(_01801_));
 sky130_fd_sc_hd__buf_1 _10378_ (.A(_05476_),
    .X(_05490_));
 sky130_fd_sc_hd__buf_1 _10379_ (.A(_05122_),
    .X(_05491_));
 sky130_fd_sc_hd__buf_1 _10380_ (.A(_05479_),
    .X(_05492_));
 sky130_fd_sc_hd__a22o_1 _10381_ (.A1(\r1.regblock[24][13] ),
    .A2(_05490_),
    .B1(_05491_),
    .B2(_05492_),
    .X(_02826_));
 sky130_fd_sc_hd__clkbuf_1 _10382_ (.A(_05488_),
    .X(_01800_));
 sky130_fd_sc_hd__buf_1 _10383_ (.A(_05125_),
    .X(_05493_));
 sky130_fd_sc_hd__a22o_1 _10384_ (.A1(\r1.regblock[24][12] ),
    .A2(_05490_),
    .B1(_05493_),
    .B2(_05492_),
    .X(_02825_));
 sky130_fd_sc_hd__clkbuf_2 _10385_ (.A(_05434_),
    .X(_05494_));
 sky130_fd_sc_hd__buf_1 _10386_ (.A(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__buf_1 _10387_ (.A(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__clkbuf_2 _10388_ (.A(_05496_),
    .X(_01799_));
 sky130_fd_sc_hd__buf_1 _10389_ (.A(_05128_),
    .X(_05497_));
 sky130_fd_sc_hd__a22o_1 _10390_ (.A1(\r1.regblock[24][11] ),
    .A2(_05490_),
    .B1(_05497_),
    .B2(_05492_),
    .X(_02824_));
 sky130_fd_sc_hd__clkbuf_1 _10391_ (.A(_05496_),
    .X(_01798_));
 sky130_fd_sc_hd__clkbuf_2 _10392_ (.A(_05453_),
    .X(_05498_));
 sky130_fd_sc_hd__buf_1 _10393_ (.A(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__buf_1 _10394_ (.A(_05132_),
    .X(_05500_));
 sky130_fd_sc_hd__clkbuf_2 _10395_ (.A(_05457_),
    .X(_05501_));
 sky130_fd_sc_hd__buf_1 _10396_ (.A(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__a22o_1 _10397_ (.A1(\r1.regblock[24][10] ),
    .A2(_05499_),
    .B1(_05500_),
    .B2(_05502_),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_1 _10398_ (.A(_05496_),
    .X(_01797_));
 sky130_fd_sc_hd__buf_1 _10399_ (.A(_05136_),
    .X(_05503_));
 sky130_fd_sc_hd__a22o_1 _10400_ (.A1(\r1.regblock[24][9] ),
    .A2(_05499_),
    .B1(_05503_),
    .B2(_05502_),
    .X(_02822_));
 sky130_fd_sc_hd__buf_1 _10401_ (.A(_05495_),
    .X(_05504_));
 sky130_fd_sc_hd__clkbuf_1 _10402_ (.A(_05504_),
    .X(_01796_));
 sky130_fd_sc_hd__buf_1 _10403_ (.A(_05142_),
    .X(_05505_));
 sky130_fd_sc_hd__a22o_1 _10404_ (.A1(\r1.regblock[24][8] ),
    .A2(_05499_),
    .B1(_05505_),
    .B2(_05502_),
    .X(_02821_));
 sky130_fd_sc_hd__clkbuf_1 _10405_ (.A(_05504_),
    .X(_01795_));
 sky130_fd_sc_hd__buf_1 _10406_ (.A(_05498_),
    .X(_05506_));
 sky130_fd_sc_hd__buf_1 _10407_ (.A(_05145_),
    .X(_05507_));
 sky130_fd_sc_hd__buf_1 _10408_ (.A(_05501_),
    .X(_05508_));
 sky130_fd_sc_hd__a22o_1 _10409_ (.A1(\r1.regblock[24][7] ),
    .A2(_05506_),
    .B1(_05507_),
    .B2(_05508_),
    .X(_02820_));
 sky130_fd_sc_hd__clkbuf_1 _10410_ (.A(_05504_),
    .X(_01794_));
 sky130_fd_sc_hd__buf_1 _10411_ (.A(_05148_),
    .X(_05509_));
 sky130_fd_sc_hd__a22o_1 _10412_ (.A1(\r1.regblock[24][6] ),
    .A2(_05506_),
    .B1(_05509_),
    .B2(_05508_),
    .X(_02819_));
 sky130_fd_sc_hd__buf_1 _10413_ (.A(_05495_),
    .X(_05510_));
 sky130_fd_sc_hd__clkbuf_1 _10414_ (.A(_05510_),
    .X(_01793_));
 sky130_fd_sc_hd__buf_1 _10415_ (.A(_05151_),
    .X(_05511_));
 sky130_fd_sc_hd__a22o_1 _10416_ (.A1(\r1.regblock[24][5] ),
    .A2(_05506_),
    .B1(_05511_),
    .B2(_05508_),
    .X(_02818_));
 sky130_fd_sc_hd__clkbuf_1 _10417_ (.A(_05510_),
    .X(_01792_));
 sky130_fd_sc_hd__buf_1 _10418_ (.A(_05498_),
    .X(_05512_));
 sky130_fd_sc_hd__buf_1 _10419_ (.A(_05154_),
    .X(_05513_));
 sky130_fd_sc_hd__buf_1 _10420_ (.A(_05501_),
    .X(_05514_));
 sky130_fd_sc_hd__a22o_1 _10421_ (.A1(\r1.regblock[24][4] ),
    .A2(_05512_),
    .B1(_05513_),
    .B2(_05514_),
    .X(_02817_));
 sky130_fd_sc_hd__clkbuf_1 _10422_ (.A(_05510_),
    .X(_01791_));
 sky130_fd_sc_hd__buf_1 _10423_ (.A(_05157_),
    .X(_05515_));
 sky130_fd_sc_hd__a22o_1 _10424_ (.A1(\r1.regblock[24][3] ),
    .A2(_05512_),
    .B1(_05515_),
    .B2(_05514_),
    .X(_02816_));
 sky130_fd_sc_hd__buf_2 _10425_ (.A(_05494_),
    .X(_05516_));
 sky130_fd_sc_hd__buf_1 _10426_ (.A(_05516_),
    .X(_05517_));
 sky130_fd_sc_hd__clkbuf_1 _10427_ (.A(_05517_),
    .X(_01790_));
 sky130_fd_sc_hd__buf_1 _10428_ (.A(_05160_),
    .X(_05518_));
 sky130_fd_sc_hd__a22o_1 _10429_ (.A1(\r1.regblock[24][2] ),
    .A2(_05512_),
    .B1(_05518_),
    .B2(_05514_),
    .X(_02815_));
 sky130_fd_sc_hd__clkbuf_1 _10430_ (.A(_05517_),
    .X(_01789_));
 sky130_fd_sc_hd__buf_1 _10431_ (.A(_05162_),
    .X(_05519_));
 sky130_fd_sc_hd__a22o_1 _10432_ (.A1(\r1.regblock[24][1] ),
    .A2(_05443_),
    .B1(_05519_),
    .B2(_05447_),
    .X(_02814_));
 sky130_fd_sc_hd__clkbuf_1 _10433_ (.A(_05517_),
    .X(_01788_));
 sky130_fd_sc_hd__buf_1 _10434_ (.A(_05164_),
    .X(_05520_));
 sky130_fd_sc_hd__a22o_1 _10435_ (.A1(\r1.regblock[24][0] ),
    .A2(_05443_),
    .B1(_05520_),
    .B2(_05447_),
    .X(_02813_));
 sky130_fd_sc_hd__buf_1 _10436_ (.A(_05516_),
    .X(_05521_));
 sky130_fd_sc_hd__clkbuf_1 _10437_ (.A(_05521_),
    .X(_01787_));
 sky130_fd_sc_hd__or2_2 _10438_ (.A(_05262_),
    .B(_04778_),
    .X(_05522_));
 sky130_fd_sc_hd__buf_1 _10439_ (.A(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__buf_1 _10440_ (.A(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__inv_2 _10441_ (.A(_05522_),
    .Y(_05525_));
 sky130_fd_sc_hd__buf_1 _10442_ (.A(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__buf_1 _10443_ (.A(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__a22o_1 _10444_ (.A1(\r1.regblock[11][31] ),
    .A2(_05524_),
    .B1(_05445_),
    .B2(_05527_),
    .X(_02812_));
 sky130_fd_sc_hd__clkbuf_1 _10445_ (.A(_05521_),
    .X(_01786_));
 sky130_fd_sc_hd__a22o_1 _10446_ (.A1(\r1.regblock[11][30] ),
    .A2(_05524_),
    .B1(_05449_),
    .B2(_05527_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_1 _10447_ (.A(_05521_),
    .X(_01785_));
 sky130_fd_sc_hd__a22o_1 _10448_ (.A1(\r1.regblock[11][29] ),
    .A2(_05524_),
    .B1(_05452_),
    .B2(_05527_),
    .X(_02810_));
 sky130_fd_sc_hd__buf_1 _10449_ (.A(_05516_),
    .X(_05528_));
 sky130_fd_sc_hd__clkbuf_1 _10450_ (.A(_05528_),
    .X(_01784_));
 sky130_fd_sc_hd__clkbuf_4 _10451_ (.A(_05522_),
    .X(_05529_));
 sky130_fd_sc_hd__clkbuf_2 _10452_ (.A(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__buf_1 _10453_ (.A(_05530_),
    .X(_05531_));
 sky130_fd_sc_hd__clkbuf_4 _10454_ (.A(_05525_),
    .X(_05532_));
 sky130_fd_sc_hd__clkbuf_2 _10455_ (.A(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__buf_1 _10456_ (.A(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__a22o_1 _10457_ (.A1(\r1.regblock[11][28] ),
    .A2(_05531_),
    .B1(_05456_),
    .B2(_05534_),
    .X(_02809_));
 sky130_fd_sc_hd__clkbuf_1 _10458_ (.A(_05528_),
    .X(_01783_));
 sky130_fd_sc_hd__a22o_1 _10459_ (.A1(\r1.regblock[11][27] ),
    .A2(_05531_),
    .B1(_05460_),
    .B2(_05534_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_1 _10460_ (.A(_05528_),
    .X(_01782_));
 sky130_fd_sc_hd__a22o_1 _10461_ (.A1(\r1.regblock[11][26] ),
    .A2(_05531_),
    .B1(_05462_),
    .B2(_05534_),
    .X(_02807_));
 sky130_fd_sc_hd__clkbuf_4 _10462_ (.A(_05494_),
    .X(_05535_));
 sky130_fd_sc_hd__buf_1 _10463_ (.A(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__clkbuf_1 _10464_ (.A(_05536_),
    .X(_01781_));
 sky130_fd_sc_hd__buf_1 _10465_ (.A(_05530_),
    .X(_05537_));
 sky130_fd_sc_hd__buf_1 _10466_ (.A(_05533_),
    .X(_05538_));
 sky130_fd_sc_hd__a22o_1 _10467_ (.A1(\r1.regblock[11][25] ),
    .A2(_05537_),
    .B1(_05464_),
    .B2(_05538_),
    .X(_02806_));
 sky130_fd_sc_hd__clkbuf_1 _10468_ (.A(_05536_),
    .X(_01780_));
 sky130_fd_sc_hd__a22o_1 _10469_ (.A1(\r1.regblock[11][24] ),
    .A2(_05537_),
    .B1(_05466_),
    .B2(_05538_),
    .X(_02805_));
 sky130_fd_sc_hd__clkbuf_1 _10470_ (.A(_05536_),
    .X(_01779_));
 sky130_fd_sc_hd__a22o_1 _10471_ (.A1(\r1.regblock[11][23] ),
    .A2(_05537_),
    .B1(_05468_),
    .B2(_05538_),
    .X(_02804_));
 sky130_fd_sc_hd__buf_1 _10472_ (.A(_05535_),
    .X(_05539_));
 sky130_fd_sc_hd__clkbuf_1 _10473_ (.A(_05539_),
    .X(_01778_));
 sky130_fd_sc_hd__buf_1 _10474_ (.A(_05530_),
    .X(_05540_));
 sky130_fd_sc_hd__buf_1 _10475_ (.A(_05533_),
    .X(_05541_));
 sky130_fd_sc_hd__a22o_1 _10476_ (.A1(\r1.regblock[11][22] ),
    .A2(_05540_),
    .B1(_05470_),
    .B2(_05541_),
    .X(_02803_));
 sky130_fd_sc_hd__clkbuf_1 _10477_ (.A(_05539_),
    .X(_01777_));
 sky130_fd_sc_hd__a22o_1 _10478_ (.A1(\r1.regblock[11][21] ),
    .A2(_05540_),
    .B1(_05472_),
    .B2(_05541_),
    .X(_02802_));
 sky130_fd_sc_hd__clkbuf_1 _10479_ (.A(_05539_),
    .X(_01776_));
 sky130_fd_sc_hd__a22o_1 _10480_ (.A1(\r1.regblock[11][20] ),
    .A2(_05540_),
    .B1(_05475_),
    .B2(_05541_),
    .X(_02801_));
 sky130_fd_sc_hd__buf_1 _10481_ (.A(_05535_),
    .X(_05542_));
 sky130_fd_sc_hd__clkbuf_1 _10482_ (.A(_05542_),
    .X(_01775_));
 sky130_fd_sc_hd__buf_2 _10483_ (.A(_05529_),
    .X(_05543_));
 sky130_fd_sc_hd__buf_1 _10484_ (.A(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__buf_2 _10485_ (.A(_05532_),
    .X(_05545_));
 sky130_fd_sc_hd__buf_1 _10486_ (.A(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__a22o_1 _10487_ (.A1(\r1.regblock[11][19] ),
    .A2(_05544_),
    .B1(_05478_),
    .B2(_05546_),
    .X(_02800_));
 sky130_fd_sc_hd__clkbuf_1 _10488_ (.A(_05542_),
    .X(_01774_));
 sky130_fd_sc_hd__a22o_1 _10489_ (.A1(\r1.regblock[11][18] ),
    .A2(_05544_),
    .B1(_05481_),
    .B2(_05546_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_1 _10490_ (.A(_05542_),
    .X(_01773_));
 sky130_fd_sc_hd__a22o_1 _10491_ (.A1(\r1.regblock[11][17] ),
    .A2(_05544_),
    .B1(_05483_),
    .B2(_05546_),
    .X(_02798_));
 sky130_fd_sc_hd__buf_1 _10492_ (.A(_05434_),
    .X(_05547_));
 sky130_fd_sc_hd__buf_4 _10493_ (.A(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__buf_1 _10494_ (.A(_05548_),
    .X(_05549_));
 sky130_fd_sc_hd__clkbuf_1 _10495_ (.A(_05549_),
    .X(_01772_));
 sky130_fd_sc_hd__buf_1 _10496_ (.A(_05543_),
    .X(_05550_));
 sky130_fd_sc_hd__buf_1 _10497_ (.A(_05545_),
    .X(_05551_));
 sky130_fd_sc_hd__a22o_1 _10498_ (.A1(\r1.regblock[11][16] ),
    .A2(_05550_),
    .B1(_05485_),
    .B2(_05551_),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_1 _10499_ (.A(_05549_),
    .X(_01771_));
 sky130_fd_sc_hd__a22o_1 _10500_ (.A1(\r1.regblock[11][15] ),
    .A2(_05550_),
    .B1(_05487_),
    .B2(_05551_),
    .X(_02796_));
 sky130_fd_sc_hd__clkbuf_1 _10501_ (.A(_05549_),
    .X(_01770_));
 sky130_fd_sc_hd__a22o_1 _10502_ (.A1(\r1.regblock[11][14] ),
    .A2(_05550_),
    .B1(_05489_),
    .B2(_05551_),
    .X(_02795_));
 sky130_fd_sc_hd__buf_1 _10503_ (.A(_05548_),
    .X(_05552_));
 sky130_fd_sc_hd__clkbuf_1 _10504_ (.A(_05552_),
    .X(_01769_));
 sky130_fd_sc_hd__buf_1 _10505_ (.A(_05543_),
    .X(_05553_));
 sky130_fd_sc_hd__buf_1 _10506_ (.A(_05545_),
    .X(_05554_));
 sky130_fd_sc_hd__a22o_1 _10507_ (.A1(\r1.regblock[11][13] ),
    .A2(_05553_),
    .B1(_05491_),
    .B2(_05554_),
    .X(_02794_));
 sky130_fd_sc_hd__clkbuf_1 _10508_ (.A(_05552_),
    .X(_01768_));
 sky130_fd_sc_hd__a22o_1 _10509_ (.A1(\r1.regblock[11][12] ),
    .A2(_05553_),
    .B1(_05493_),
    .B2(_05554_),
    .X(_02793_));
 sky130_fd_sc_hd__clkbuf_1 _10510_ (.A(_05552_),
    .X(_01767_));
 sky130_fd_sc_hd__a22o_1 _10511_ (.A1(\r1.regblock[11][11] ),
    .A2(_05553_),
    .B1(_05497_),
    .B2(_05554_),
    .X(_02792_));
 sky130_fd_sc_hd__buf_1 _10512_ (.A(_05548_),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_1 _10513_ (.A(_05555_),
    .X(_01766_));
 sky130_fd_sc_hd__clkbuf_2 _10514_ (.A(_05529_),
    .X(_05556_));
 sky130_fd_sc_hd__buf_1 _10515_ (.A(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__clkbuf_2 _10516_ (.A(_05532_),
    .X(_05558_));
 sky130_fd_sc_hd__buf_1 _10517_ (.A(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__a22o_1 _10518_ (.A1(\r1.regblock[11][10] ),
    .A2(_05557_),
    .B1(_05500_),
    .B2(_05559_),
    .X(_02791_));
 sky130_fd_sc_hd__clkbuf_1 _10519_ (.A(_05555_),
    .X(_01765_));
 sky130_fd_sc_hd__a22o_1 _10520_ (.A1(\r1.regblock[11][9] ),
    .A2(_05557_),
    .B1(_05503_),
    .B2(_05559_),
    .X(_02790_));
 sky130_fd_sc_hd__clkbuf_1 _10521_ (.A(_05555_),
    .X(_01764_));
 sky130_fd_sc_hd__a22o_1 _10522_ (.A1(\r1.regblock[11][8] ),
    .A2(_05557_),
    .B1(_05505_),
    .B2(_05559_),
    .X(_02789_));
 sky130_fd_sc_hd__buf_2 _10523_ (.A(_05547_),
    .X(_05560_));
 sky130_fd_sc_hd__buf_1 _10524_ (.A(_05560_),
    .X(_05561_));
 sky130_fd_sc_hd__clkbuf_1 _10525_ (.A(_05561_),
    .X(_01763_));
 sky130_fd_sc_hd__buf_1 _10526_ (.A(_05556_),
    .X(_05562_));
 sky130_fd_sc_hd__buf_1 _10527_ (.A(_05558_),
    .X(_05563_));
 sky130_fd_sc_hd__a22o_1 _10528_ (.A1(\r1.regblock[11][7] ),
    .A2(_05562_),
    .B1(_05507_),
    .B2(_05563_),
    .X(_02788_));
 sky130_fd_sc_hd__clkbuf_1 _10529_ (.A(_05561_),
    .X(_01762_));
 sky130_fd_sc_hd__a22o_1 _10530_ (.A1(\r1.regblock[11][6] ),
    .A2(_05562_),
    .B1(_05509_),
    .B2(_05563_),
    .X(_02787_));
 sky130_fd_sc_hd__clkbuf_1 _10531_ (.A(_05561_),
    .X(_01761_));
 sky130_fd_sc_hd__a22o_1 _10532_ (.A1(\r1.regblock[11][5] ),
    .A2(_05562_),
    .B1(_05511_),
    .B2(_05563_),
    .X(_02786_));
 sky130_fd_sc_hd__buf_1 _10533_ (.A(_05560_),
    .X(_05564_));
 sky130_fd_sc_hd__clkbuf_1 _10534_ (.A(_05564_),
    .X(_01760_));
 sky130_fd_sc_hd__buf_1 _10535_ (.A(_05556_),
    .X(_05565_));
 sky130_fd_sc_hd__buf_1 _10536_ (.A(_05558_),
    .X(_05566_));
 sky130_fd_sc_hd__a22o_1 _10537_ (.A1(\r1.regblock[11][4] ),
    .A2(_05565_),
    .B1(_05513_),
    .B2(_05566_),
    .X(_02785_));
 sky130_fd_sc_hd__clkbuf_1 _10538_ (.A(_05564_),
    .X(_01759_));
 sky130_fd_sc_hd__a22o_1 _10539_ (.A1(\r1.regblock[11][3] ),
    .A2(_05565_),
    .B1(_05515_),
    .B2(_05566_),
    .X(_02784_));
 sky130_fd_sc_hd__clkbuf_1 _10540_ (.A(_05564_),
    .X(_01758_));
 sky130_fd_sc_hd__a22o_1 _10541_ (.A1(\r1.regblock[11][2] ),
    .A2(_05565_),
    .B1(_05518_),
    .B2(_05566_),
    .X(_02783_));
 sky130_fd_sc_hd__buf_1 _10542_ (.A(_05560_),
    .X(_05567_));
 sky130_fd_sc_hd__clkbuf_1 _10543_ (.A(_05567_),
    .X(_01757_));
 sky130_fd_sc_hd__a22o_1 _10544_ (.A1(\r1.regblock[11][1] ),
    .A2(_05523_),
    .B1(_05519_),
    .B2(_05526_),
    .X(_02782_));
 sky130_fd_sc_hd__clkbuf_1 _10545_ (.A(_05567_),
    .X(_01756_));
 sky130_fd_sc_hd__a22o_1 _10546_ (.A1(\r1.regblock[11][0] ),
    .A2(_05523_),
    .B1(_05520_),
    .B2(_05526_),
    .X(_02781_));
 sky130_fd_sc_hd__clkbuf_1 _10547_ (.A(_05567_),
    .X(_01755_));
 sky130_fd_sc_hd__or2_2 _10548_ (.A(_05054_),
    .B(_04777_),
    .X(_05568_));
 sky130_fd_sc_hd__buf_1 _10549_ (.A(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__buf_1 _10550_ (.A(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__inv_2 _10551_ (.A(_05568_),
    .Y(_05571_));
 sky130_fd_sc_hd__buf_1 _10552_ (.A(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__buf_1 _10553_ (.A(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__a22o_1 _10554_ (.A1(\r1.regblock[10][31] ),
    .A2(_05570_),
    .B1(_05445_),
    .B2(_05573_),
    .X(_02780_));
 sky130_fd_sc_hd__clkbuf_2 _10555_ (.A(_05547_),
    .X(_05574_));
 sky130_fd_sc_hd__buf_1 _10556_ (.A(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__clkbuf_1 _10557_ (.A(_05575_),
    .X(_01754_));
 sky130_fd_sc_hd__a22o_1 _10558_ (.A1(\r1.regblock[10][30] ),
    .A2(_05570_),
    .B1(_05449_),
    .B2(_05573_),
    .X(_02779_));
 sky130_fd_sc_hd__clkbuf_1 _10559_ (.A(_05575_),
    .X(_01753_));
 sky130_fd_sc_hd__a22o_1 _10560_ (.A1(\r1.regblock[10][29] ),
    .A2(_05570_),
    .B1(_05452_),
    .B2(_05573_),
    .X(_02778_));
 sky130_fd_sc_hd__clkbuf_1 _10561_ (.A(_05575_),
    .X(_01752_));
 sky130_fd_sc_hd__clkbuf_4 _10562_ (.A(_05568_),
    .X(_05576_));
 sky130_fd_sc_hd__clkbuf_2 _10563_ (.A(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__buf_1 _10564_ (.A(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__clkbuf_4 _10565_ (.A(_05571_),
    .X(_05579_));
 sky130_fd_sc_hd__clkbuf_2 _10566_ (.A(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__buf_1 _10567_ (.A(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__a22o_1 _10568_ (.A1(\r1.regblock[10][28] ),
    .A2(_05578_),
    .B1(_05456_),
    .B2(_05581_),
    .X(_02777_));
 sky130_fd_sc_hd__buf_1 _10569_ (.A(_05574_),
    .X(_05582_));
 sky130_fd_sc_hd__clkbuf_1 _10570_ (.A(_05582_),
    .X(_01751_));
 sky130_fd_sc_hd__a22o_1 _10571_ (.A1(\r1.regblock[10][27] ),
    .A2(_05578_),
    .B1(_05460_),
    .B2(_05581_),
    .X(_02776_));
 sky130_fd_sc_hd__clkbuf_1 _10572_ (.A(_05582_),
    .X(_01750_));
 sky130_fd_sc_hd__a22o_1 _10573_ (.A1(\r1.regblock[10][26] ),
    .A2(_05578_),
    .B1(_05462_),
    .B2(_05581_),
    .X(_02775_));
 sky130_fd_sc_hd__clkbuf_1 _10574_ (.A(_05582_),
    .X(_01749_));
 sky130_fd_sc_hd__buf_1 _10575_ (.A(_05577_),
    .X(_05583_));
 sky130_fd_sc_hd__buf_1 _10576_ (.A(_05580_),
    .X(_05584_));
 sky130_fd_sc_hd__a22o_1 _10577_ (.A1(\r1.regblock[10][25] ),
    .A2(_05583_),
    .B1(_05464_),
    .B2(_05584_),
    .X(_02774_));
 sky130_fd_sc_hd__buf_1 _10578_ (.A(_05574_),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_1 _10579_ (.A(_05585_),
    .X(_01748_));
 sky130_fd_sc_hd__a22o_1 _10580_ (.A1(\r1.regblock[10][24] ),
    .A2(_05583_),
    .B1(_05466_),
    .B2(_05584_),
    .X(_02773_));
 sky130_fd_sc_hd__clkbuf_1 _10581_ (.A(_05585_),
    .X(_01747_));
 sky130_fd_sc_hd__a22o_1 _10582_ (.A1(\r1.regblock[10][23] ),
    .A2(_05583_),
    .B1(_05468_),
    .B2(_05584_),
    .X(_02772_));
 sky130_fd_sc_hd__buf_1 _10583_ (.A(_05585_),
    .X(_01746_));
 sky130_fd_sc_hd__buf_1 _10584_ (.A(_05577_),
    .X(_05586_));
 sky130_fd_sc_hd__buf_1 _10585_ (.A(_05580_),
    .X(_05587_));
 sky130_fd_sc_hd__a22o_1 _10586_ (.A1(\r1.regblock[10][22] ),
    .A2(_05586_),
    .B1(_05470_),
    .B2(_05587_),
    .X(_02771_));
 sky130_fd_sc_hd__buf_1 _10587_ (.A(_05433_),
    .X(_05588_));
 sky130_fd_sc_hd__clkbuf_2 _10588_ (.A(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__clkbuf_2 _10589_ (.A(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__buf_2 _10590_ (.A(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__clkbuf_1 _10591_ (.A(_05591_),
    .X(_01745_));
 sky130_fd_sc_hd__a22o_1 _10592_ (.A1(\r1.regblock[10][21] ),
    .A2(_05586_),
    .B1(_05472_),
    .B2(_05587_),
    .X(_02770_));
 sky130_fd_sc_hd__clkbuf_1 _10593_ (.A(_05591_),
    .X(_01744_));
 sky130_fd_sc_hd__a22o_1 _10594_ (.A1(\r1.regblock[10][20] ),
    .A2(_05586_),
    .B1(_05475_),
    .B2(_05587_),
    .X(_02769_));
 sky130_fd_sc_hd__clkbuf_1 _10595_ (.A(_05591_),
    .X(_01743_));
 sky130_fd_sc_hd__clkbuf_2 _10596_ (.A(_05576_),
    .X(_05592_));
 sky130_fd_sc_hd__buf_1 _10597_ (.A(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__clkbuf_2 _10598_ (.A(_05579_),
    .X(_05594_));
 sky130_fd_sc_hd__buf_1 _10599_ (.A(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__a22o_1 _10600_ (.A1(\r1.regblock[10][19] ),
    .A2(_05593_),
    .B1(_05478_),
    .B2(_05595_),
    .X(_02768_));
 sky130_fd_sc_hd__buf_1 _10601_ (.A(_05590_),
    .X(_05596_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(_05596_),
    .X(_01742_));
 sky130_fd_sc_hd__a22o_1 _10603_ (.A1(\r1.regblock[10][18] ),
    .A2(_05593_),
    .B1(_05481_),
    .B2(_05595_),
    .X(_02767_));
 sky130_fd_sc_hd__clkbuf_1 _10604_ (.A(_05596_),
    .X(_01741_));
 sky130_fd_sc_hd__a22o_1 _10605_ (.A1(\r1.regblock[10][17] ),
    .A2(_05593_),
    .B1(_05483_),
    .B2(_05595_),
    .X(_02766_));
 sky130_fd_sc_hd__clkbuf_1 _10606_ (.A(_05596_),
    .X(_01740_));
 sky130_fd_sc_hd__buf_1 _10607_ (.A(_05592_),
    .X(_05597_));
 sky130_fd_sc_hd__buf_1 _10608_ (.A(_05594_),
    .X(_05598_));
 sky130_fd_sc_hd__a22o_1 _10609_ (.A1(\r1.regblock[10][16] ),
    .A2(_05597_),
    .B1(_05485_),
    .B2(_05598_),
    .X(_02765_));
 sky130_fd_sc_hd__buf_1 _10610_ (.A(_05590_),
    .X(_05599_));
 sky130_fd_sc_hd__clkbuf_1 _10611_ (.A(_05599_),
    .X(_01739_));
 sky130_fd_sc_hd__a22o_1 _10612_ (.A1(\r1.regblock[10][15] ),
    .A2(_05597_),
    .B1(_05487_),
    .B2(_05598_),
    .X(_02764_));
 sky130_fd_sc_hd__clkbuf_1 _10613_ (.A(_05599_),
    .X(_01738_));
 sky130_fd_sc_hd__a22o_1 _10614_ (.A1(\r1.regblock[10][14] ),
    .A2(_05597_),
    .B1(_05489_),
    .B2(_05598_),
    .X(_02763_));
 sky130_fd_sc_hd__clkbuf_1 _10615_ (.A(_05599_),
    .X(_01737_));
 sky130_fd_sc_hd__buf_1 _10616_ (.A(_05592_),
    .X(_05600_));
 sky130_fd_sc_hd__buf_1 _10617_ (.A(_05594_),
    .X(_05601_));
 sky130_fd_sc_hd__a22o_1 _10618_ (.A1(\r1.regblock[10][13] ),
    .A2(_05600_),
    .B1(_05491_),
    .B2(_05601_),
    .X(_02762_));
 sky130_fd_sc_hd__clkbuf_2 _10619_ (.A(_05589_),
    .X(_05602_));
 sky130_fd_sc_hd__buf_2 _10620_ (.A(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__clkbuf_1 _10621_ (.A(_05603_),
    .X(_01736_));
 sky130_fd_sc_hd__a22o_1 _10622_ (.A1(\r1.regblock[10][12] ),
    .A2(_05600_),
    .B1(_05493_),
    .B2(_05601_),
    .X(_02761_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(_05603_),
    .X(_01735_));
 sky130_fd_sc_hd__a22o_1 _10624_ (.A1(\r1.regblock[10][11] ),
    .A2(_05600_),
    .B1(_05497_),
    .B2(_05601_),
    .X(_02760_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(_05603_),
    .X(_01734_));
 sky130_fd_sc_hd__clkbuf_2 _10626_ (.A(_05576_),
    .X(_05604_));
 sky130_fd_sc_hd__buf_1 _10627_ (.A(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__clkbuf_2 _10628_ (.A(_05579_),
    .X(_05606_));
 sky130_fd_sc_hd__buf_1 _10629_ (.A(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__a22o_1 _10630_ (.A1(\r1.regblock[10][10] ),
    .A2(_05605_),
    .B1(_05500_),
    .B2(_05607_),
    .X(_02759_));
 sky130_fd_sc_hd__buf_1 _10631_ (.A(_05602_),
    .X(_05608_));
 sky130_fd_sc_hd__clkbuf_1 _10632_ (.A(_05608_),
    .X(_01733_));
 sky130_fd_sc_hd__a22o_1 _10633_ (.A1(\r1.regblock[10][9] ),
    .A2(_05605_),
    .B1(_05503_),
    .B2(_05607_),
    .X(_02758_));
 sky130_fd_sc_hd__clkbuf_1 _10634_ (.A(_05608_),
    .X(_01732_));
 sky130_fd_sc_hd__a22o_1 _10635_ (.A1(\r1.regblock[10][8] ),
    .A2(_05605_),
    .B1(_05505_),
    .B2(_05607_),
    .X(_02757_));
 sky130_fd_sc_hd__clkbuf_1 _10636_ (.A(_05608_),
    .X(_01731_));
 sky130_fd_sc_hd__buf_1 _10637_ (.A(_05604_),
    .X(_05609_));
 sky130_fd_sc_hd__buf_1 _10638_ (.A(_05606_),
    .X(_05610_));
 sky130_fd_sc_hd__a22o_1 _10639_ (.A1(\r1.regblock[10][7] ),
    .A2(_05609_),
    .B1(_05507_),
    .B2(_05610_),
    .X(_02756_));
 sky130_fd_sc_hd__buf_1 _10640_ (.A(_05602_),
    .X(_05611_));
 sky130_fd_sc_hd__clkbuf_1 _10641_ (.A(_05611_),
    .X(_01730_));
 sky130_fd_sc_hd__a22o_1 _10642_ (.A1(\r1.regblock[10][6] ),
    .A2(_05609_),
    .B1(_05509_),
    .B2(_05610_),
    .X(_02755_));
 sky130_fd_sc_hd__clkbuf_1 _10643_ (.A(_05611_),
    .X(_01729_));
 sky130_fd_sc_hd__a22o_1 _10644_ (.A1(\r1.regblock[10][5] ),
    .A2(_05609_),
    .B1(_05511_),
    .B2(_05610_),
    .X(_02754_));
 sky130_fd_sc_hd__clkbuf_1 _10645_ (.A(_05611_),
    .X(_01728_));
 sky130_fd_sc_hd__buf_1 _10646_ (.A(_05604_),
    .X(_05612_));
 sky130_fd_sc_hd__buf_1 _10647_ (.A(_05606_),
    .X(_05613_));
 sky130_fd_sc_hd__a22o_1 _10648_ (.A1(\r1.regblock[10][4] ),
    .A2(_05612_),
    .B1(_05513_),
    .B2(_05613_),
    .X(_02753_));
 sky130_fd_sc_hd__buf_1 _10649_ (.A(_05589_),
    .X(_05614_));
 sky130_fd_sc_hd__clkbuf_2 _10650_ (.A(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__clkbuf_1 _10651_ (.A(_05615_),
    .X(_01727_));
 sky130_fd_sc_hd__a22o_1 _10652_ (.A1(\r1.regblock[10][3] ),
    .A2(_05612_),
    .B1(_05515_),
    .B2(_05613_),
    .X(_02752_));
 sky130_fd_sc_hd__clkbuf_1 _10653_ (.A(_05615_),
    .X(_01726_));
 sky130_fd_sc_hd__a22o_1 _10654_ (.A1(\r1.regblock[10][2] ),
    .A2(_05612_),
    .B1(_05518_),
    .B2(_05613_),
    .X(_02751_));
 sky130_fd_sc_hd__clkbuf_1 _10655_ (.A(_05615_),
    .X(_01725_));
 sky130_fd_sc_hd__a22o_1 _10656_ (.A1(\r1.regblock[10][1] ),
    .A2(_05569_),
    .B1(_05519_),
    .B2(_05572_),
    .X(_02750_));
 sky130_fd_sc_hd__buf_1 _10657_ (.A(_05614_),
    .X(_05616_));
 sky130_fd_sc_hd__clkbuf_1 _10658_ (.A(_05616_),
    .X(_01724_));
 sky130_fd_sc_hd__a22o_1 _10659_ (.A1(\r1.regblock[10][0] ),
    .A2(_05569_),
    .B1(_05520_),
    .B2(_05572_),
    .X(_02749_));
 sky130_fd_sc_hd__clkbuf_1 _10660_ (.A(_05616_),
    .X(_01723_));
 sky130_fd_sc_hd__or2_2 _10661_ (.A(_04449_),
    .B(_04643_),
    .X(_05617_));
 sky130_fd_sc_hd__buf_1 _10662_ (.A(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__buf_1 _10663_ (.A(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__buf_1 _10664_ (.A(_04453_),
    .X(_05620_));
 sky130_fd_sc_hd__clkbuf_2 _10665_ (.A(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__inv_2 _10666_ (.A(_05617_),
    .Y(_05622_));
 sky130_fd_sc_hd__buf_1 _10667_ (.A(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__buf_1 _10668_ (.A(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__a22o_1 _10669_ (.A1(\r1.regblock[6][31] ),
    .A2(_05619_),
    .B1(_05621_),
    .B2(_05624_),
    .X(_02748_));
 sky130_fd_sc_hd__clkbuf_1 _10670_ (.A(_05616_),
    .X(_01722_));
 sky130_fd_sc_hd__buf_1 _10671_ (.A(_04459_),
    .X(_05625_));
 sky130_fd_sc_hd__buf_1 _10672_ (.A(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__a22o_1 _10673_ (.A1(\r1.regblock[6][30] ),
    .A2(_05619_),
    .B1(_05626_),
    .B2(_05624_),
    .X(_02747_));
 sky130_fd_sc_hd__buf_2 _10674_ (.A(_05614_),
    .X(_05627_));
 sky130_fd_sc_hd__clkbuf_1 _10675_ (.A(_05627_),
    .X(_01721_));
 sky130_fd_sc_hd__buf_1 _10676_ (.A(_04463_),
    .X(_05628_));
 sky130_fd_sc_hd__buf_1 _10677_ (.A(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__a22o_1 _10678_ (.A1(\r1.regblock[6][29] ),
    .A2(_05619_),
    .B1(_05629_),
    .B2(_05624_),
    .X(_02746_));
 sky130_fd_sc_hd__clkbuf_1 _10679_ (.A(_05627_),
    .X(_01720_));
 sky130_fd_sc_hd__buf_4 _10680_ (.A(_05617_),
    .X(_05630_));
 sky130_fd_sc_hd__clkbuf_2 _10681_ (.A(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__buf_1 _10682_ (.A(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__clkbuf_2 _10683_ (.A(_04469_),
    .X(_05633_));
 sky130_fd_sc_hd__buf_1 _10684_ (.A(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__buf_4 _10685_ (.A(_05622_),
    .X(_05635_));
 sky130_fd_sc_hd__clkbuf_2 _10686_ (.A(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__buf_1 _10687_ (.A(_05636_),
    .X(_05637_));
 sky130_fd_sc_hd__a22o_1 _10688_ (.A1(\r1.regblock[6][28] ),
    .A2(_05632_),
    .B1(_05634_),
    .B2(_05637_),
    .X(_02745_));
 sky130_fd_sc_hd__clkbuf_1 _10689_ (.A(_05627_),
    .X(_01719_));
 sky130_fd_sc_hd__clkbuf_2 _10690_ (.A(_04475_),
    .X(_05638_));
 sky130_fd_sc_hd__buf_1 _10691_ (.A(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__a22o_1 _10692_ (.A1(\r1.regblock[6][27] ),
    .A2(_05632_),
    .B1(_05639_),
    .B2(_05637_),
    .X(_02744_));
 sky130_fd_sc_hd__clkbuf_4 _10693_ (.A(_05588_),
    .X(_05640_));
 sky130_fd_sc_hd__buf_1 _10694_ (.A(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__buf_1 _10695_ (.A(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__clkbuf_1 _10696_ (.A(_05642_),
    .X(_01718_));
 sky130_fd_sc_hd__clkbuf_2 _10697_ (.A(_04480_),
    .X(_05643_));
 sky130_fd_sc_hd__buf_1 _10698_ (.A(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__a22o_1 _10699_ (.A1(\r1.regblock[6][26] ),
    .A2(_05632_),
    .B1(_05644_),
    .B2(_05637_),
    .X(_02743_));
 sky130_fd_sc_hd__clkbuf_1 _10700_ (.A(_05642_),
    .X(_01717_));
 sky130_fd_sc_hd__buf_1 _10701_ (.A(_05631_),
    .X(_05645_));
 sky130_fd_sc_hd__clkbuf_2 _10702_ (.A(_04484_),
    .X(_05646_));
 sky130_fd_sc_hd__buf_1 _10703_ (.A(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__buf_1 _10704_ (.A(_05636_),
    .X(_05648_));
 sky130_fd_sc_hd__a22o_1 _10705_ (.A1(\r1.regblock[6][25] ),
    .A2(_05645_),
    .B1(_05647_),
    .B2(_05648_),
    .X(_02742_));
 sky130_fd_sc_hd__clkbuf_1 _10706_ (.A(_05642_),
    .X(_01716_));
 sky130_fd_sc_hd__buf_1 _10707_ (.A(_04488_),
    .X(_05649_));
 sky130_fd_sc_hd__buf_1 _10708_ (.A(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__a22o_1 _10709_ (.A1(\r1.regblock[6][24] ),
    .A2(_05645_),
    .B1(_05650_),
    .B2(_05648_),
    .X(_02741_));
 sky130_fd_sc_hd__buf_1 _10710_ (.A(_05641_),
    .X(_05651_));
 sky130_fd_sc_hd__clkbuf_1 _10711_ (.A(_05651_),
    .X(_01715_));
 sky130_fd_sc_hd__buf_1 _10712_ (.A(_04492_),
    .X(_05652_));
 sky130_fd_sc_hd__buf_1 _10713_ (.A(_05652_),
    .X(_05653_));
 sky130_fd_sc_hd__a22o_1 _10714_ (.A1(\r1.regblock[6][23] ),
    .A2(_05645_),
    .B1(_05653_),
    .B2(_05648_),
    .X(_02740_));
 sky130_fd_sc_hd__clkbuf_1 _10715_ (.A(_05651_),
    .X(_01714_));
 sky130_fd_sc_hd__buf_1 _10716_ (.A(_05631_),
    .X(_05654_));
 sky130_fd_sc_hd__buf_1 _10717_ (.A(_04496_),
    .X(_05655_));
 sky130_fd_sc_hd__buf_1 _10718_ (.A(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__buf_1 _10719_ (.A(_05636_),
    .X(_05657_));
 sky130_fd_sc_hd__a22o_1 _10720_ (.A1(\r1.regblock[6][22] ),
    .A2(_05654_),
    .B1(_05656_),
    .B2(_05657_),
    .X(_02739_));
 sky130_fd_sc_hd__clkbuf_1 _10721_ (.A(_05651_),
    .X(_01713_));
 sky130_fd_sc_hd__buf_1 _10722_ (.A(_04500_),
    .X(_05658_));
 sky130_fd_sc_hd__buf_1 _10723_ (.A(_05658_),
    .X(_05659_));
 sky130_fd_sc_hd__a22o_1 _10724_ (.A1(\r1.regblock[6][21] ),
    .A2(_05654_),
    .B1(_05659_),
    .B2(_05657_),
    .X(_02738_));
 sky130_fd_sc_hd__clkbuf_4 _10725_ (.A(_05641_),
    .X(_05660_));
 sky130_fd_sc_hd__clkbuf_1 _10726_ (.A(_05660_),
    .X(_01712_));
 sky130_fd_sc_hd__clkbuf_2 _10727_ (.A(_04504_),
    .X(_05661_));
 sky130_fd_sc_hd__buf_1 _10728_ (.A(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__a22o_1 _10729_ (.A1(\r1.regblock[6][20] ),
    .A2(_05654_),
    .B1(_05662_),
    .B2(_05657_),
    .X(_02737_));
 sky130_fd_sc_hd__clkbuf_1 _10730_ (.A(_05660_),
    .X(_01711_));
 sky130_fd_sc_hd__buf_1 _10731_ (.A(_05630_),
    .X(_05663_));
 sky130_fd_sc_hd__buf_1 _10732_ (.A(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__clkbuf_2 _10733_ (.A(_04509_),
    .X(_05665_));
 sky130_fd_sc_hd__buf_1 _10734_ (.A(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__buf_1 _10735_ (.A(_05635_),
    .X(_05667_));
 sky130_fd_sc_hd__buf_1 _10736_ (.A(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__a22o_1 _10737_ (.A1(\r1.regblock[6][19] ),
    .A2(_05664_),
    .B1(_05666_),
    .B2(_05668_),
    .X(_02736_));
 sky130_fd_sc_hd__clkbuf_1 _10738_ (.A(_05660_),
    .X(_01710_));
 sky130_fd_sc_hd__clkbuf_2 _10739_ (.A(_04514_),
    .X(_05669_));
 sky130_fd_sc_hd__buf_1 _10740_ (.A(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__a22o_1 _10741_ (.A1(\r1.regblock[6][18] ),
    .A2(_05664_),
    .B1(_05670_),
    .B2(_05668_),
    .X(_02735_));
 sky130_fd_sc_hd__buf_1 _10742_ (.A(_05640_),
    .X(_05671_));
 sky130_fd_sc_hd__buf_1 _10743_ (.A(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__clkbuf_1 _10744_ (.A(_05672_),
    .X(_01709_));
 sky130_fd_sc_hd__clkbuf_2 _10745_ (.A(_04520_),
    .X(_05673_));
 sky130_fd_sc_hd__buf_1 _10746_ (.A(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__a22o_1 _10747_ (.A1(\r1.regblock[6][17] ),
    .A2(_05664_),
    .B1(_05674_),
    .B2(_05668_),
    .X(_02734_));
 sky130_fd_sc_hd__clkbuf_1 _10748_ (.A(_05672_),
    .X(_01708_));
 sky130_fd_sc_hd__buf_1 _10749_ (.A(_05663_),
    .X(_05675_));
 sky130_fd_sc_hd__buf_2 _10750_ (.A(_04524_),
    .X(_05676_));
 sky130_fd_sc_hd__buf_1 _10751_ (.A(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__buf_1 _10752_ (.A(_05667_),
    .X(_05678_));
 sky130_fd_sc_hd__a22o_1 _10753_ (.A1(\r1.regblock[6][16] ),
    .A2(_05675_),
    .B1(_05677_),
    .B2(_05678_),
    .X(_02733_));
 sky130_fd_sc_hd__clkbuf_1 _10754_ (.A(_05672_),
    .X(_01707_));
 sky130_fd_sc_hd__clkbuf_2 _10755_ (.A(_04528_),
    .X(_05679_));
 sky130_fd_sc_hd__clkbuf_2 _10756_ (.A(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__a22o_1 _10757_ (.A1(\r1.regblock[6][15] ),
    .A2(_05675_),
    .B1(_05680_),
    .B2(_05678_),
    .X(_02732_));
 sky130_fd_sc_hd__buf_1 _10758_ (.A(_05671_),
    .X(_05681_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(_05681_),
    .X(_01706_));
 sky130_fd_sc_hd__clkbuf_2 _10760_ (.A(_04532_),
    .X(_05682_));
 sky130_fd_sc_hd__clkbuf_2 _10761_ (.A(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__a22o_1 _10762_ (.A1(\r1.regblock[6][14] ),
    .A2(_05675_),
    .B1(_05683_),
    .B2(_05678_),
    .X(_02731_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(_05681_),
    .X(_01705_));
 sky130_fd_sc_hd__buf_1 _10764_ (.A(_05663_),
    .X(_05684_));
 sky130_fd_sc_hd__buf_2 _10765_ (.A(_04536_),
    .X(_05685_));
 sky130_fd_sc_hd__buf_1 _10766_ (.A(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__buf_1 _10767_ (.A(_05667_),
    .X(_05687_));
 sky130_fd_sc_hd__a22o_1 _10768_ (.A1(\r1.regblock[6][13] ),
    .A2(_05684_),
    .B1(_05686_),
    .B2(_05687_),
    .X(_02730_));
 sky130_fd_sc_hd__clkbuf_1 _10769_ (.A(_05681_),
    .X(_01704_));
 sky130_fd_sc_hd__buf_2 _10770_ (.A(_04540_),
    .X(_05688_));
 sky130_fd_sc_hd__buf_1 _10771_ (.A(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__a22o_1 _10772_ (.A1(\r1.regblock[6][12] ),
    .A2(_05684_),
    .B1(_05689_),
    .B2(_05687_),
    .X(_02729_));
 sky130_fd_sc_hd__buf_2 _10773_ (.A(_05671_),
    .X(_05690_));
 sky130_fd_sc_hd__clkbuf_1 _10774_ (.A(_05690_),
    .X(_01703_));
 sky130_fd_sc_hd__clkbuf_2 _10775_ (.A(_04544_),
    .X(_05691_));
 sky130_fd_sc_hd__buf_1 _10776_ (.A(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__a22o_1 _10777_ (.A1(\r1.regblock[6][11] ),
    .A2(_05684_),
    .B1(_05692_),
    .B2(_05687_),
    .X(_02728_));
 sky130_fd_sc_hd__clkbuf_1 _10778_ (.A(_05690_),
    .X(_01702_));
 sky130_fd_sc_hd__buf_1 _10779_ (.A(_05630_),
    .X(_05693_));
 sky130_fd_sc_hd__buf_1 _10780_ (.A(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__buf_1 _10781_ (.A(_04549_),
    .X(_05695_));
 sky130_fd_sc_hd__clkbuf_2 _10782_ (.A(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__buf_1 _10783_ (.A(_05635_),
    .X(_05697_));
 sky130_fd_sc_hd__buf_1 _10784_ (.A(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__a22o_1 _10785_ (.A1(\r1.regblock[6][10] ),
    .A2(_05694_),
    .B1(_05696_),
    .B2(_05698_),
    .X(_02727_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(_05690_),
    .X(_01701_));
 sky130_fd_sc_hd__clkbuf_2 _10787_ (.A(_04554_),
    .X(_05699_));
 sky130_fd_sc_hd__buf_1 _10788_ (.A(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__a22o_1 _10789_ (.A1(\r1.regblock[6][9] ),
    .A2(_05694_),
    .B1(_05700_),
    .B2(_05698_),
    .X(_02726_));
 sky130_fd_sc_hd__buf_1 _10790_ (.A(_05640_),
    .X(_05701_));
 sky130_fd_sc_hd__buf_1 _10791_ (.A(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(_05702_),
    .X(_01700_));
 sky130_fd_sc_hd__clkbuf_2 _10793_ (.A(_04559_),
    .X(_05703_));
 sky130_fd_sc_hd__buf_1 _10794_ (.A(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__a22o_1 _10795_ (.A1(\r1.regblock[6][8] ),
    .A2(_05694_),
    .B1(_05704_),
    .B2(_05698_),
    .X(_02725_));
 sky130_fd_sc_hd__clkbuf_1 _10796_ (.A(_05702_),
    .X(_01699_));
 sky130_fd_sc_hd__buf_1 _10797_ (.A(_05693_),
    .X(_05705_));
 sky130_fd_sc_hd__clkbuf_2 _10798_ (.A(_04563_),
    .X(_05706_));
 sky130_fd_sc_hd__buf_1 _10799_ (.A(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__buf_1 _10800_ (.A(_05697_),
    .X(_05708_));
 sky130_fd_sc_hd__a22o_1 _10801_ (.A1(\r1.regblock[6][7] ),
    .A2(_05705_),
    .B1(_05707_),
    .B2(_05708_),
    .X(_02724_));
 sky130_fd_sc_hd__clkbuf_1 _10802_ (.A(_05702_),
    .X(_01698_));
 sky130_fd_sc_hd__clkbuf_2 _10803_ (.A(_04567_),
    .X(_05709_));
 sky130_fd_sc_hd__buf_1 _10804_ (.A(_05709_),
    .X(_05710_));
 sky130_fd_sc_hd__a22o_1 _10805_ (.A1(\r1.regblock[6][6] ),
    .A2(_05705_),
    .B1(_05710_),
    .B2(_05708_),
    .X(_02723_));
 sky130_fd_sc_hd__buf_1 _10806_ (.A(_05701_),
    .X(_05711_));
 sky130_fd_sc_hd__clkbuf_1 _10807_ (.A(_05711_),
    .X(_01697_));
 sky130_fd_sc_hd__clkbuf_2 _10808_ (.A(_04571_),
    .X(_05712_));
 sky130_fd_sc_hd__buf_1 _10809_ (.A(_05712_),
    .X(_05713_));
 sky130_fd_sc_hd__a22o_1 _10810_ (.A1(\r1.regblock[6][5] ),
    .A2(_05705_),
    .B1(_05713_),
    .B2(_05708_),
    .X(_02722_));
 sky130_fd_sc_hd__clkbuf_1 _10811_ (.A(_05711_),
    .X(_01696_));
 sky130_fd_sc_hd__buf_1 _10812_ (.A(_05693_),
    .X(_05714_));
 sky130_fd_sc_hd__clkbuf_2 _10813_ (.A(_04575_),
    .X(_05715_));
 sky130_fd_sc_hd__buf_1 _10814_ (.A(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__buf_1 _10815_ (.A(_05697_),
    .X(_05717_));
 sky130_fd_sc_hd__a22o_1 _10816_ (.A1(\r1.regblock[6][4] ),
    .A2(_05714_),
    .B1(_05716_),
    .B2(_05717_),
    .X(_02721_));
 sky130_fd_sc_hd__clkbuf_1 _10817_ (.A(_05711_),
    .X(_01695_));
 sky130_fd_sc_hd__clkbuf_2 _10818_ (.A(_04579_),
    .X(_05718_));
 sky130_fd_sc_hd__buf_1 _10819_ (.A(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__a22o_1 _10820_ (.A1(\r1.regblock[6][3] ),
    .A2(_05714_),
    .B1(_05719_),
    .B2(_05717_),
    .X(_02720_));
 sky130_fd_sc_hd__buf_2 _10821_ (.A(_05701_),
    .X(_05720_));
 sky130_fd_sc_hd__clkbuf_1 _10822_ (.A(_05720_),
    .X(_01694_));
 sky130_fd_sc_hd__clkbuf_2 _10823_ (.A(_04583_),
    .X(_05721_));
 sky130_fd_sc_hd__buf_1 _10824_ (.A(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__a22o_1 _10825_ (.A1(\r1.regblock[6][2] ),
    .A2(_05714_),
    .B1(_05722_),
    .B2(_05717_),
    .X(_02719_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(_05720_),
    .X(_01693_));
 sky130_fd_sc_hd__buf_1 _10827_ (.A(_04586_),
    .X(_05723_));
 sky130_fd_sc_hd__buf_1 _10828_ (.A(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__a22o_1 _10829_ (.A1(\r1.regblock[6][1] ),
    .A2(_05618_),
    .B1(_05724_),
    .B2(_05623_),
    .X(_02718_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(_05720_),
    .X(_01692_));
 sky130_fd_sc_hd__buf_1 _10831_ (.A(_04589_),
    .X(_05725_));
 sky130_fd_sc_hd__buf_1 _10832_ (.A(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__a22o_1 _10833_ (.A1(\r1.regblock[6][0] ),
    .A2(_05618_),
    .B1(_05726_),
    .B2(_05623_),
    .X(_02717_));
 sky130_fd_sc_hd__buf_1 _10834_ (.A(_05588_),
    .X(_05727_));
 sky130_fd_sc_hd__buf_2 _10835_ (.A(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__buf_1 _10836_ (.A(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__clkbuf_1 _10837_ (.A(_05729_),
    .X(_01691_));
 sky130_fd_sc_hd__or2_2 _10838_ (.A(_05262_),
    .B(_04642_),
    .X(_05730_));
 sky130_fd_sc_hd__buf_1 _10839_ (.A(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__buf_1 _10840_ (.A(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__inv_2 _10841_ (.A(_05730_),
    .Y(_05733_));
 sky130_fd_sc_hd__buf_1 _10842_ (.A(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__buf_1 _10843_ (.A(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__a22o_1 _10844_ (.A1(\r1.regblock[7][31] ),
    .A2(_05732_),
    .B1(_05621_),
    .B2(_05735_),
    .X(_02716_));
 sky130_fd_sc_hd__clkbuf_1 _10845_ (.A(_05729_),
    .X(_01690_));
 sky130_fd_sc_hd__a22o_1 _10846_ (.A1(\r1.regblock[7][30] ),
    .A2(_05732_),
    .B1(_05626_),
    .B2(_05735_),
    .X(_02715_));
 sky130_fd_sc_hd__clkbuf_1 _10847_ (.A(_05729_),
    .X(_01689_));
 sky130_fd_sc_hd__a22o_1 _10848_ (.A1(\r1.regblock[7][29] ),
    .A2(_05732_),
    .B1(_05629_),
    .B2(_05735_),
    .X(_02714_));
 sky130_fd_sc_hd__buf_1 _10849_ (.A(_05728_),
    .X(_05736_));
 sky130_fd_sc_hd__clkbuf_1 _10850_ (.A(_05736_),
    .X(_01688_));
 sky130_fd_sc_hd__buf_4 _10851_ (.A(_05730_),
    .X(_05737_));
 sky130_fd_sc_hd__clkbuf_2 _10852_ (.A(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__buf_1 _10853_ (.A(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__buf_4 _10854_ (.A(_05733_),
    .X(_05740_));
 sky130_fd_sc_hd__clkbuf_2 _10855_ (.A(_05740_),
    .X(_05741_));
 sky130_fd_sc_hd__buf_1 _10856_ (.A(_05741_),
    .X(_05742_));
 sky130_fd_sc_hd__a22o_1 _10857_ (.A1(\r1.regblock[7][28] ),
    .A2(_05739_),
    .B1(_05634_),
    .B2(_05742_),
    .X(_02713_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(_05736_),
    .X(_01687_));
 sky130_fd_sc_hd__a22o_1 _10859_ (.A1(\r1.regblock[7][27] ),
    .A2(_05739_),
    .B1(_05639_),
    .B2(_05742_),
    .X(_02712_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_05736_),
    .X(_01686_));
 sky130_fd_sc_hd__a22o_1 _10861_ (.A1(\r1.regblock[7][26] ),
    .A2(_05739_),
    .B1(_05644_),
    .B2(_05742_),
    .X(_02711_));
 sky130_fd_sc_hd__buf_1 _10862_ (.A(_05728_),
    .X(_05743_));
 sky130_fd_sc_hd__clkbuf_1 _10863_ (.A(_05743_),
    .X(_01685_));
 sky130_fd_sc_hd__buf_1 _10864_ (.A(_05738_),
    .X(_05744_));
 sky130_fd_sc_hd__buf_1 _10865_ (.A(_05741_),
    .X(_05745_));
 sky130_fd_sc_hd__a22o_1 _10866_ (.A1(\r1.regblock[7][25] ),
    .A2(_05744_),
    .B1(_05647_),
    .B2(_05745_),
    .X(_02710_));
 sky130_fd_sc_hd__clkbuf_1 _10867_ (.A(_05743_),
    .X(_01684_));
 sky130_fd_sc_hd__a22o_1 _10868_ (.A1(\r1.regblock[7][24] ),
    .A2(_05744_),
    .B1(_05650_),
    .B2(_05745_),
    .X(_02709_));
 sky130_fd_sc_hd__clkbuf_1 _10869_ (.A(_05743_),
    .X(_01683_));
 sky130_fd_sc_hd__a22o_1 _10870_ (.A1(\r1.regblock[7][23] ),
    .A2(_05744_),
    .B1(_05653_),
    .B2(_05745_),
    .X(_02708_));
 sky130_fd_sc_hd__clkbuf_4 _10871_ (.A(_05727_),
    .X(_05746_));
 sky130_fd_sc_hd__buf_1 _10872_ (.A(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__clkbuf_1 _10873_ (.A(_05747_),
    .X(_01682_));
 sky130_fd_sc_hd__buf_1 _10874_ (.A(_05738_),
    .X(_05748_));
 sky130_fd_sc_hd__buf_1 _10875_ (.A(_05741_),
    .X(_05749_));
 sky130_fd_sc_hd__a22o_1 _10876_ (.A1(\r1.regblock[7][22] ),
    .A2(_05748_),
    .B1(_05656_),
    .B2(_05749_),
    .X(_02707_));
 sky130_fd_sc_hd__clkbuf_1 _10877_ (.A(_05747_),
    .X(_01681_));
 sky130_fd_sc_hd__a22o_1 _10878_ (.A1(\r1.regblock[7][21] ),
    .A2(_05748_),
    .B1(_05659_),
    .B2(_05749_),
    .X(_02706_));
 sky130_fd_sc_hd__clkbuf_1 _10879_ (.A(_05747_),
    .X(_01680_));
 sky130_fd_sc_hd__a22o_1 _10880_ (.A1(\r1.regblock[7][20] ),
    .A2(_05748_),
    .B1(_05662_),
    .B2(_05749_),
    .X(_02705_));
 sky130_fd_sc_hd__buf_1 _10881_ (.A(_05746_),
    .X(_05750_));
 sky130_fd_sc_hd__clkbuf_1 _10882_ (.A(_05750_),
    .X(_01679_));
 sky130_fd_sc_hd__buf_1 _10883_ (.A(_05737_),
    .X(_05751_));
 sky130_fd_sc_hd__buf_1 _10884_ (.A(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__buf_1 _10885_ (.A(_05740_),
    .X(_05753_));
 sky130_fd_sc_hd__buf_1 _10886_ (.A(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__a22o_1 _10887_ (.A1(\r1.regblock[7][19] ),
    .A2(_05752_),
    .B1(_05666_),
    .B2(_05754_),
    .X(_02704_));
 sky130_fd_sc_hd__clkbuf_1 _10888_ (.A(_05750_),
    .X(_01678_));
 sky130_fd_sc_hd__a22o_1 _10889_ (.A1(\r1.regblock[7][18] ),
    .A2(_05752_),
    .B1(_05670_),
    .B2(_05754_),
    .X(_02703_));
 sky130_fd_sc_hd__clkbuf_1 _10890_ (.A(_05750_),
    .X(_01677_));
 sky130_fd_sc_hd__a22o_1 _10891_ (.A1(\r1.regblock[7][17] ),
    .A2(_05752_),
    .B1(_05674_),
    .B2(_05754_),
    .X(_02702_));
 sky130_fd_sc_hd__buf_1 _10892_ (.A(_05746_),
    .X(_05755_));
 sky130_fd_sc_hd__clkbuf_1 _10893_ (.A(_05755_),
    .X(_01676_));
 sky130_fd_sc_hd__buf_1 _10894_ (.A(_05751_),
    .X(_05756_));
 sky130_fd_sc_hd__buf_1 _10895_ (.A(_05753_),
    .X(_05757_));
 sky130_fd_sc_hd__a22o_1 _10896_ (.A1(\r1.regblock[7][16] ),
    .A2(_05756_),
    .B1(_05677_),
    .B2(_05757_),
    .X(_02701_));
 sky130_fd_sc_hd__clkbuf_1 _10897_ (.A(_05755_),
    .X(_01675_));
 sky130_fd_sc_hd__a22o_1 _10898_ (.A1(\r1.regblock[7][15] ),
    .A2(_05756_),
    .B1(_05680_),
    .B2(_05757_),
    .X(_02700_));
 sky130_fd_sc_hd__clkbuf_1 _10899_ (.A(_05755_),
    .X(_01674_));
 sky130_fd_sc_hd__a22o_1 _10900_ (.A1(\r1.regblock[7][14] ),
    .A2(_05756_),
    .B1(_05683_),
    .B2(_05757_),
    .X(_02699_));
 sky130_fd_sc_hd__buf_4 _10901_ (.A(_05727_),
    .X(_05758_));
 sky130_fd_sc_hd__buf_1 _10902_ (.A(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__clkbuf_1 _10903_ (.A(_05759_),
    .X(_01673_));
 sky130_fd_sc_hd__buf_1 _10904_ (.A(_05751_),
    .X(_05760_));
 sky130_fd_sc_hd__buf_1 _10905_ (.A(_05753_),
    .X(_05761_));
 sky130_fd_sc_hd__a22o_1 _10906_ (.A1(\r1.regblock[7][13] ),
    .A2(_05760_),
    .B1(_05686_),
    .B2(_05761_),
    .X(_02698_));
 sky130_fd_sc_hd__clkbuf_1 _10907_ (.A(_05759_),
    .X(_01672_));
 sky130_fd_sc_hd__a22o_1 _10908_ (.A1(\r1.regblock[7][12] ),
    .A2(_05760_),
    .B1(_05689_),
    .B2(_05761_),
    .X(_02697_));
 sky130_fd_sc_hd__clkbuf_1 _10909_ (.A(_05759_),
    .X(_01671_));
 sky130_fd_sc_hd__a22o_1 _10910_ (.A1(\r1.regblock[7][11] ),
    .A2(_05760_),
    .B1(_05692_),
    .B2(_05761_),
    .X(_02696_));
 sky130_fd_sc_hd__buf_1 _10911_ (.A(_05758_),
    .X(_05762_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(_05762_),
    .X(_01670_));
 sky130_fd_sc_hd__buf_1 _10913_ (.A(_05737_),
    .X(_05763_));
 sky130_fd_sc_hd__buf_1 _10914_ (.A(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__buf_1 _10915_ (.A(_05740_),
    .X(_05765_));
 sky130_fd_sc_hd__buf_1 _10916_ (.A(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__a22o_1 _10917_ (.A1(\r1.regblock[7][10] ),
    .A2(_05764_),
    .B1(_05696_),
    .B2(_05766_),
    .X(_02695_));
 sky130_fd_sc_hd__clkbuf_1 _10918_ (.A(_05762_),
    .X(_01669_));
 sky130_fd_sc_hd__a22o_1 _10919_ (.A1(\r1.regblock[7][9] ),
    .A2(_05764_),
    .B1(_05700_),
    .B2(_05766_),
    .X(_02694_));
 sky130_fd_sc_hd__clkbuf_1 _10920_ (.A(_05762_),
    .X(_01668_));
 sky130_fd_sc_hd__a22o_1 _10921_ (.A1(\r1.regblock[7][8] ),
    .A2(_05764_),
    .B1(_05704_),
    .B2(_05766_),
    .X(_02693_));
 sky130_fd_sc_hd__buf_1 _10922_ (.A(_05758_),
    .X(_05767_));
 sky130_fd_sc_hd__clkbuf_1 _10923_ (.A(_05767_),
    .X(_01667_));
 sky130_fd_sc_hd__buf_1 _10924_ (.A(_05763_),
    .X(_05768_));
 sky130_fd_sc_hd__buf_1 _10925_ (.A(_05765_),
    .X(_05769_));
 sky130_fd_sc_hd__a22o_1 _10926_ (.A1(\r1.regblock[7][7] ),
    .A2(_05768_),
    .B1(_05707_),
    .B2(_05769_),
    .X(_02692_));
 sky130_fd_sc_hd__clkbuf_1 _10927_ (.A(_05767_),
    .X(_01666_));
 sky130_fd_sc_hd__a22o_1 _10928_ (.A1(\r1.regblock[7][6] ),
    .A2(_05768_),
    .B1(_05710_),
    .B2(_05769_),
    .X(_02691_));
 sky130_fd_sc_hd__clkbuf_1 _10929_ (.A(_05767_),
    .X(_01665_));
 sky130_fd_sc_hd__a22o_1 _10930_ (.A1(\r1.regblock[7][5] ),
    .A2(_05768_),
    .B1(_05713_),
    .B2(_05769_),
    .X(_02690_));
 sky130_fd_sc_hd__buf_1 _10931_ (.A(_05433_),
    .X(_05770_));
 sky130_fd_sc_hd__buf_2 _10932_ (.A(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__buf_2 _10933_ (.A(_05771_),
    .X(_05772_));
 sky130_fd_sc_hd__buf_1 _10934_ (.A(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__clkbuf_1 _10935_ (.A(_05773_),
    .X(_01664_));
 sky130_fd_sc_hd__buf_1 _10936_ (.A(_05763_),
    .X(_05774_));
 sky130_fd_sc_hd__buf_1 _10937_ (.A(_05765_),
    .X(_05775_));
 sky130_fd_sc_hd__a22o_1 _10938_ (.A1(\r1.regblock[7][4] ),
    .A2(_05774_),
    .B1(_05716_),
    .B2(_05775_),
    .X(_02689_));
 sky130_fd_sc_hd__clkbuf_1 _10939_ (.A(_05773_),
    .X(_01663_));
 sky130_fd_sc_hd__a22o_1 _10940_ (.A1(\r1.regblock[7][3] ),
    .A2(_05774_),
    .B1(_05719_),
    .B2(_05775_),
    .X(_02688_));
 sky130_fd_sc_hd__clkbuf_1 _10941_ (.A(_05773_),
    .X(_01662_));
 sky130_fd_sc_hd__a22o_1 _10942_ (.A1(\r1.regblock[7][2] ),
    .A2(_05774_),
    .B1(_05722_),
    .B2(_05775_),
    .X(_02687_));
 sky130_fd_sc_hd__buf_1 _10943_ (.A(_05772_),
    .X(_05776_));
 sky130_fd_sc_hd__clkbuf_1 _10944_ (.A(_05776_),
    .X(_01661_));
 sky130_fd_sc_hd__a22o_1 _10945_ (.A1(\r1.regblock[7][1] ),
    .A2(_05731_),
    .B1(_05724_),
    .B2(_05734_),
    .X(_02686_));
 sky130_fd_sc_hd__clkbuf_1 _10946_ (.A(_05776_),
    .X(_01660_));
 sky130_fd_sc_hd__a22o_1 _10947_ (.A1(\r1.regblock[7][0] ),
    .A2(_05731_),
    .B1(_05726_),
    .B2(_05734_),
    .X(_02685_));
 sky130_fd_sc_hd__clkbuf_1 _10948_ (.A(_05776_),
    .X(_01659_));
 sky130_fd_sc_hd__or2_2 _10949_ (.A(_04643_),
    .B(_04775_),
    .X(_05777_));
 sky130_fd_sc_hd__buf_1 _10950_ (.A(_05777_),
    .X(_05778_));
 sky130_fd_sc_hd__buf_1 _10951_ (.A(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__inv_2 _10952_ (.A(_05777_),
    .Y(_05780_));
 sky130_fd_sc_hd__buf_1 _10953_ (.A(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__buf_1 _10954_ (.A(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__a22o_1 _10955_ (.A1(\r1.regblock[4][31] ),
    .A2(_05779_),
    .B1(_05621_),
    .B2(_05782_),
    .X(_02684_));
 sky130_fd_sc_hd__clkbuf_2 _10956_ (.A(_05772_),
    .X(_05783_));
 sky130_fd_sc_hd__clkbuf_1 _10957_ (.A(_05783_),
    .X(_01658_));
 sky130_fd_sc_hd__a22o_1 _10958_ (.A1(\r1.regblock[4][30] ),
    .A2(_05779_),
    .B1(_05626_),
    .B2(_05782_),
    .X(_02683_));
 sky130_fd_sc_hd__clkbuf_1 _10959_ (.A(_05783_),
    .X(_01657_));
 sky130_fd_sc_hd__a22o_1 _10960_ (.A1(\r1.regblock[4][29] ),
    .A2(_05779_),
    .B1(_05629_),
    .B2(_05782_),
    .X(_02682_));
 sky130_fd_sc_hd__clkbuf_1 _10961_ (.A(_05783_),
    .X(_01656_));
 sky130_fd_sc_hd__buf_4 _10962_ (.A(_05777_),
    .X(_05784_));
 sky130_fd_sc_hd__clkbuf_2 _10963_ (.A(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__buf_1 _10964_ (.A(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__buf_4 _10965_ (.A(_05780_),
    .X(_05787_));
 sky130_fd_sc_hd__clkbuf_2 _10966_ (.A(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__buf_1 _10967_ (.A(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__a22o_1 _10968_ (.A1(\r1.regblock[4][28] ),
    .A2(_05786_),
    .B1(_05634_),
    .B2(_05789_),
    .X(_02681_));
 sky130_fd_sc_hd__clkbuf_2 _10969_ (.A(_05771_),
    .X(_05790_));
 sky130_fd_sc_hd__buf_1 _10970_ (.A(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__clkbuf_1 _10971_ (.A(_05791_),
    .X(_01655_));
 sky130_fd_sc_hd__a22o_1 _10972_ (.A1(\r1.regblock[4][27] ),
    .A2(_05786_),
    .B1(_05639_),
    .B2(_05789_),
    .X(_02680_));
 sky130_fd_sc_hd__clkbuf_1 _10973_ (.A(_05791_),
    .X(_01654_));
 sky130_fd_sc_hd__a22o_1 _10974_ (.A1(\r1.regblock[4][26] ),
    .A2(_05786_),
    .B1(_05644_),
    .B2(_05789_),
    .X(_02679_));
 sky130_fd_sc_hd__clkbuf_1 _10975_ (.A(_05791_),
    .X(_01653_));
 sky130_fd_sc_hd__buf_1 _10976_ (.A(_05785_),
    .X(_05792_));
 sky130_fd_sc_hd__buf_1 _10977_ (.A(_05788_),
    .X(_05793_));
 sky130_fd_sc_hd__a22o_1 _10978_ (.A1(\r1.regblock[4][25] ),
    .A2(_05792_),
    .B1(_05647_),
    .B2(_05793_),
    .X(_02678_));
 sky130_fd_sc_hd__buf_1 _10979_ (.A(_05790_),
    .X(_05794_));
 sky130_fd_sc_hd__clkbuf_1 _10980_ (.A(_05794_),
    .X(_01652_));
 sky130_fd_sc_hd__a22o_1 _10981_ (.A1(\r1.regblock[4][24] ),
    .A2(_05792_),
    .B1(_05650_),
    .B2(_05793_),
    .X(_02677_));
 sky130_fd_sc_hd__clkbuf_1 _10982_ (.A(_05794_),
    .X(_01651_));
 sky130_fd_sc_hd__a22o_1 _10983_ (.A1(\r1.regblock[4][23] ),
    .A2(_05792_),
    .B1(_05653_),
    .B2(_05793_),
    .X(_02676_));
 sky130_fd_sc_hd__clkbuf_1 _10984_ (.A(_05794_),
    .X(_01650_));
 sky130_fd_sc_hd__buf_1 _10985_ (.A(_05785_),
    .X(_05795_));
 sky130_fd_sc_hd__buf_1 _10986_ (.A(_05788_),
    .X(_05796_));
 sky130_fd_sc_hd__a22o_1 _10987_ (.A1(\r1.regblock[4][22] ),
    .A2(_05795_),
    .B1(_05656_),
    .B2(_05796_),
    .X(_02675_));
 sky130_fd_sc_hd__buf_1 _10988_ (.A(_05790_),
    .X(_05797_));
 sky130_fd_sc_hd__clkbuf_1 _10989_ (.A(_05797_),
    .X(_01649_));
 sky130_fd_sc_hd__a22o_1 _10990_ (.A1(\r1.regblock[4][21] ),
    .A2(_05795_),
    .B1(_05659_),
    .B2(_05796_),
    .X(_02674_));
 sky130_fd_sc_hd__clkbuf_1 _10991_ (.A(_05797_),
    .X(_01648_));
 sky130_fd_sc_hd__a22o_1 _10992_ (.A1(\r1.regblock[4][20] ),
    .A2(_05795_),
    .B1(_05662_),
    .B2(_05796_),
    .X(_02673_));
 sky130_fd_sc_hd__buf_2 _10993_ (.A(_05797_),
    .X(_01647_));
 sky130_fd_sc_hd__buf_1 _10994_ (.A(_05784_),
    .X(_05798_));
 sky130_fd_sc_hd__buf_1 _10995_ (.A(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__buf_1 _10996_ (.A(_05787_),
    .X(_05800_));
 sky130_fd_sc_hd__buf_1 _10997_ (.A(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__a22o_1 _10998_ (.A1(\r1.regblock[4][19] ),
    .A2(_05799_),
    .B1(_05666_),
    .B2(_05801_),
    .X(_02672_));
 sky130_fd_sc_hd__clkbuf_2 _10999_ (.A(_05771_),
    .X(_05802_));
 sky130_fd_sc_hd__buf_1 _11000_ (.A(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__clkbuf_1 _11001_ (.A(_05803_),
    .X(_01646_));
 sky130_fd_sc_hd__a22o_1 _11002_ (.A1(\r1.regblock[4][18] ),
    .A2(_05799_),
    .B1(_05670_),
    .B2(_05801_),
    .X(_02671_));
 sky130_fd_sc_hd__clkbuf_1 _11003_ (.A(_05803_),
    .X(_01645_));
 sky130_fd_sc_hd__a22o_1 _11004_ (.A1(\r1.regblock[4][17] ),
    .A2(_05799_),
    .B1(_05674_),
    .B2(_05801_),
    .X(_02670_));
 sky130_fd_sc_hd__clkbuf_1 _11005_ (.A(_05803_),
    .X(_01644_));
 sky130_fd_sc_hd__buf_1 _11006_ (.A(_05798_),
    .X(_05804_));
 sky130_fd_sc_hd__buf_1 _11007_ (.A(_05800_),
    .X(_05805_));
 sky130_fd_sc_hd__a22o_1 _11008_ (.A1(\r1.regblock[4][16] ),
    .A2(_05804_),
    .B1(_05677_),
    .B2(_05805_),
    .X(_02669_));
 sky130_fd_sc_hd__buf_1 _11009_ (.A(_05802_),
    .X(_05806_));
 sky130_fd_sc_hd__clkbuf_1 _11010_ (.A(_05806_),
    .X(_01643_));
 sky130_fd_sc_hd__a22o_1 _11011_ (.A1(\r1.regblock[4][15] ),
    .A2(_05804_),
    .B1(_05680_),
    .B2(_05805_),
    .X(_02668_));
 sky130_fd_sc_hd__clkbuf_1 _11012_ (.A(_05806_),
    .X(_01642_));
 sky130_fd_sc_hd__a22o_1 _11013_ (.A1(\r1.regblock[4][14] ),
    .A2(_05804_),
    .B1(_05683_),
    .B2(_05805_),
    .X(_02667_));
 sky130_fd_sc_hd__clkbuf_1 _11014_ (.A(_05806_),
    .X(_01641_));
 sky130_fd_sc_hd__buf_1 _11015_ (.A(_05798_),
    .X(_05807_));
 sky130_fd_sc_hd__buf_1 _11016_ (.A(_05800_),
    .X(_05808_));
 sky130_fd_sc_hd__a22o_1 _11017_ (.A1(\r1.regblock[4][13] ),
    .A2(_05807_),
    .B1(_05686_),
    .B2(_05808_),
    .X(_02666_));
 sky130_fd_sc_hd__buf_1 _11018_ (.A(_05802_),
    .X(_05809_));
 sky130_fd_sc_hd__clkbuf_1 _11019_ (.A(_05809_),
    .X(_01640_));
 sky130_fd_sc_hd__a22o_1 _11020_ (.A1(\r1.regblock[4][12] ),
    .A2(_05807_),
    .B1(_05689_),
    .B2(_05808_),
    .X(_02665_));
 sky130_fd_sc_hd__clkbuf_1 _11021_ (.A(_05809_),
    .X(_01639_));
 sky130_fd_sc_hd__a22o_1 _11022_ (.A1(\r1.regblock[4][11] ),
    .A2(_05807_),
    .B1(_05692_),
    .B2(_05808_),
    .X(_02664_));
 sky130_fd_sc_hd__clkbuf_2 _11023_ (.A(_05809_),
    .X(_01638_));
 sky130_fd_sc_hd__buf_1 _11024_ (.A(_05784_),
    .X(_05810_));
 sky130_fd_sc_hd__buf_1 _11025_ (.A(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__buf_1 _11026_ (.A(_05787_),
    .X(_05812_));
 sky130_fd_sc_hd__buf_1 _11027_ (.A(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__a22o_1 _11028_ (.A1(\r1.regblock[4][10] ),
    .A2(_05811_),
    .B1(_05696_),
    .B2(_05813_),
    .X(_02663_));
 sky130_fd_sc_hd__clkbuf_2 _11029_ (.A(_05770_),
    .X(_05814_));
 sky130_fd_sc_hd__clkbuf_2 _11030_ (.A(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__buf_1 _11031_ (.A(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__clkbuf_1 _11032_ (.A(_05816_),
    .X(_01637_));
 sky130_fd_sc_hd__a22o_1 _11033_ (.A1(\r1.regblock[4][9] ),
    .A2(_05811_),
    .B1(_05700_),
    .B2(_05813_),
    .X(_02662_));
 sky130_fd_sc_hd__clkbuf_1 _11034_ (.A(_05816_),
    .X(_01636_));
 sky130_fd_sc_hd__a22o_1 _11035_ (.A1(\r1.regblock[4][8] ),
    .A2(_05811_),
    .B1(_05704_),
    .B2(_05813_),
    .X(_02661_));
 sky130_fd_sc_hd__clkbuf_1 _11036_ (.A(_05816_),
    .X(_01635_));
 sky130_fd_sc_hd__buf_1 _11037_ (.A(_05810_),
    .X(_05817_));
 sky130_fd_sc_hd__buf_1 _11038_ (.A(_05812_),
    .X(_05818_));
 sky130_fd_sc_hd__a22o_1 _11039_ (.A1(\r1.regblock[4][7] ),
    .A2(_05817_),
    .B1(_05707_),
    .B2(_05818_),
    .X(_02660_));
 sky130_fd_sc_hd__buf_1 _11040_ (.A(_05815_),
    .X(_05819_));
 sky130_fd_sc_hd__clkbuf_1 _11041_ (.A(_05819_),
    .X(_01634_));
 sky130_fd_sc_hd__a22o_1 _11042_ (.A1(\r1.regblock[4][6] ),
    .A2(_05817_),
    .B1(_05710_),
    .B2(_05818_),
    .X(_02659_));
 sky130_fd_sc_hd__clkbuf_1 _11043_ (.A(_05819_),
    .X(_01633_));
 sky130_fd_sc_hd__a22o_1 _11044_ (.A1(\r1.regblock[4][5] ),
    .A2(_05817_),
    .B1(_05713_),
    .B2(_05818_),
    .X(_02658_));
 sky130_fd_sc_hd__clkbuf_1 _11045_ (.A(_05819_),
    .X(_01632_));
 sky130_fd_sc_hd__buf_1 _11046_ (.A(_05810_),
    .X(_05820_));
 sky130_fd_sc_hd__buf_1 _11047_ (.A(_05812_),
    .X(_05821_));
 sky130_fd_sc_hd__a22o_1 _11048_ (.A1(\r1.regblock[4][4] ),
    .A2(_05820_),
    .B1(_05716_),
    .B2(_05821_),
    .X(_02657_));
 sky130_fd_sc_hd__buf_1 _11049_ (.A(_05815_),
    .X(_05822_));
 sky130_fd_sc_hd__clkbuf_1 _11050_ (.A(_05822_),
    .X(_01631_));
 sky130_fd_sc_hd__a22o_1 _11051_ (.A1(\r1.regblock[4][3] ),
    .A2(_05820_),
    .B1(_05719_),
    .B2(_05821_),
    .X(_02656_));
 sky130_fd_sc_hd__clkbuf_1 _11052_ (.A(_05822_),
    .X(_01630_));
 sky130_fd_sc_hd__a22o_1 _11053_ (.A1(\r1.regblock[4][2] ),
    .A2(_05820_),
    .B1(_05722_),
    .B2(_05821_),
    .X(_02655_));
 sky130_fd_sc_hd__buf_1 _11054_ (.A(_05822_),
    .X(_01629_));
 sky130_fd_sc_hd__a22o_1 _11055_ (.A1(\r1.regblock[4][1] ),
    .A2(_05778_),
    .B1(_05724_),
    .B2(_05781_),
    .X(_02654_));
 sky130_fd_sc_hd__clkbuf_2 _11056_ (.A(_05814_),
    .X(_05823_));
 sky130_fd_sc_hd__clkbuf_2 _11057_ (.A(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__clkbuf_1 _11058_ (.A(_05824_),
    .X(_01628_));
 sky130_fd_sc_hd__a22o_1 _11059_ (.A1(\r1.regblock[4][0] ),
    .A2(_05778_),
    .B1(_05726_),
    .B2(_05781_),
    .X(_02653_));
 sky130_fd_sc_hd__clkbuf_1 _11060_ (.A(_05824_),
    .X(_01627_));
 sky130_fd_sc_hd__clkbuf_1 _11061_ (.A(_04342_),
    .X(_05825_));
 sky130_fd_sc_hd__or2_2 _11062_ (.A(_05825_),
    .B(_04775_),
    .X(_05826_));
 sky130_fd_sc_hd__buf_1 _11063_ (.A(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__buf_1 _11064_ (.A(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__buf_1 _11065_ (.A(_05620_),
    .X(_05829_));
 sky130_fd_sc_hd__inv_2 _11066_ (.A(_05826_),
    .Y(_05830_));
 sky130_fd_sc_hd__buf_1 _11067_ (.A(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__buf_1 _11068_ (.A(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__a22o_1 _11069_ (.A1(\r1.regblock[16][31] ),
    .A2(_05828_),
    .B1(_05829_),
    .B2(_05832_),
    .X(_02652_));
 sky130_fd_sc_hd__clkbuf_1 _11070_ (.A(_05824_),
    .X(_01626_));
 sky130_fd_sc_hd__buf_1 _11071_ (.A(_05625_),
    .X(_05833_));
 sky130_fd_sc_hd__a22o_1 _11072_ (.A1(\r1.regblock[16][30] ),
    .A2(_05828_),
    .B1(_05833_),
    .B2(_05832_),
    .X(_02651_));
 sky130_fd_sc_hd__clkbuf_2 _11073_ (.A(_05823_),
    .X(_05834_));
 sky130_fd_sc_hd__clkbuf_1 _11074_ (.A(_05834_),
    .X(_01625_));
 sky130_fd_sc_hd__buf_1 _11075_ (.A(_05628_),
    .X(_05835_));
 sky130_fd_sc_hd__a22o_1 _11076_ (.A1(\r1.regblock[16][29] ),
    .A2(_05828_),
    .B1(_05835_),
    .B2(_05832_),
    .X(_02650_));
 sky130_fd_sc_hd__clkbuf_1 _11077_ (.A(_05834_),
    .X(_01624_));
 sky130_fd_sc_hd__buf_2 _11078_ (.A(_05826_),
    .X(_05836_));
 sky130_fd_sc_hd__buf_2 _11079_ (.A(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__buf_1 _11080_ (.A(_05837_),
    .X(_05838_));
 sky130_fd_sc_hd__buf_1 _11081_ (.A(_05633_),
    .X(_05839_));
 sky130_fd_sc_hd__buf_2 _11082_ (.A(_05830_),
    .X(_05840_));
 sky130_fd_sc_hd__buf_2 _11083_ (.A(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__buf_1 _11084_ (.A(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__a22o_1 _11085_ (.A1(\r1.regblock[16][28] ),
    .A2(_05838_),
    .B1(_05839_),
    .B2(_05842_),
    .X(_02649_));
 sky130_fd_sc_hd__clkbuf_1 _11086_ (.A(_05834_),
    .X(_01623_));
 sky130_fd_sc_hd__buf_1 _11087_ (.A(_05638_),
    .X(_05843_));
 sky130_fd_sc_hd__a22o_1 _11088_ (.A1(\r1.regblock[16][27] ),
    .A2(_05838_),
    .B1(_05843_),
    .B2(_05842_),
    .X(_02648_));
 sky130_fd_sc_hd__buf_1 _11089_ (.A(_05823_),
    .X(_05844_));
 sky130_fd_sc_hd__clkbuf_1 _11090_ (.A(_05844_),
    .X(_01622_));
 sky130_fd_sc_hd__buf_1 _11091_ (.A(_05643_),
    .X(_05845_));
 sky130_fd_sc_hd__a22o_1 _11092_ (.A1(\r1.regblock[16][26] ),
    .A2(_05838_),
    .B1(_05845_),
    .B2(_05842_),
    .X(_02647_));
 sky130_fd_sc_hd__clkbuf_1 _11093_ (.A(_05844_),
    .X(_01621_));
 sky130_fd_sc_hd__buf_1 _11094_ (.A(_05837_),
    .X(_05846_));
 sky130_fd_sc_hd__buf_1 _11095_ (.A(_05646_),
    .X(_05847_));
 sky130_fd_sc_hd__buf_1 _11096_ (.A(_05841_),
    .X(_05848_));
 sky130_fd_sc_hd__a22o_1 _11097_ (.A1(\r1.regblock[16][25] ),
    .A2(_05846_),
    .B1(_05847_),
    .B2(_05848_),
    .X(_02646_));
 sky130_fd_sc_hd__clkbuf_1 _11098_ (.A(_05844_),
    .X(_01620_));
 sky130_fd_sc_hd__buf_1 _11099_ (.A(_05649_),
    .X(_05849_));
 sky130_fd_sc_hd__a22o_1 _11100_ (.A1(\r1.regblock[16][24] ),
    .A2(_05846_),
    .B1(_05849_),
    .B2(_05848_),
    .X(_02645_));
 sky130_fd_sc_hd__buf_1 _11101_ (.A(_05814_),
    .X(_05850_));
 sky130_fd_sc_hd__clkbuf_2 _11102_ (.A(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__buf_1 _11103_ (.A(_05851_),
    .X(_01619_));
 sky130_fd_sc_hd__buf_1 _11104_ (.A(_05652_),
    .X(_05852_));
 sky130_fd_sc_hd__a22o_1 _11105_ (.A1(\r1.regblock[16][23] ),
    .A2(_05846_),
    .B1(_05852_),
    .B2(_05848_),
    .X(_02644_));
 sky130_fd_sc_hd__clkbuf_1 _11106_ (.A(_05851_),
    .X(_01618_));
 sky130_fd_sc_hd__buf_1 _11107_ (.A(_05837_),
    .X(_05853_));
 sky130_fd_sc_hd__buf_1 _11108_ (.A(_05655_),
    .X(_05854_));
 sky130_fd_sc_hd__buf_1 _11109_ (.A(_05841_),
    .X(_05855_));
 sky130_fd_sc_hd__a22o_1 _11110_ (.A1(\r1.regblock[16][22] ),
    .A2(_05853_),
    .B1(_05854_),
    .B2(_05855_),
    .X(_02643_));
 sky130_fd_sc_hd__clkbuf_1 _11111_ (.A(_05851_),
    .X(_01617_));
 sky130_fd_sc_hd__buf_1 _11112_ (.A(_05658_),
    .X(_05856_));
 sky130_fd_sc_hd__a22o_1 _11113_ (.A1(\r1.regblock[16][21] ),
    .A2(_05853_),
    .B1(_05856_),
    .B2(_05855_),
    .X(_02642_));
 sky130_fd_sc_hd__buf_1 _11114_ (.A(_05850_),
    .X(_05857_));
 sky130_fd_sc_hd__clkbuf_2 _11115_ (.A(_05857_),
    .X(_01616_));
 sky130_fd_sc_hd__buf_1 _11116_ (.A(_05661_),
    .X(_05858_));
 sky130_fd_sc_hd__a22o_1 _11117_ (.A1(\r1.regblock[16][20] ),
    .A2(_05853_),
    .B1(_05858_),
    .B2(_05855_),
    .X(_02641_));
 sky130_fd_sc_hd__clkbuf_1 _11118_ (.A(_05857_),
    .X(_01615_));
 sky130_fd_sc_hd__buf_2 _11119_ (.A(_05836_),
    .X(_05859_));
 sky130_fd_sc_hd__buf_1 _11120_ (.A(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__buf_1 _11121_ (.A(_05665_),
    .X(_05861_));
 sky130_fd_sc_hd__buf_2 _11122_ (.A(_05840_),
    .X(_05862_));
 sky130_fd_sc_hd__buf_1 _11123_ (.A(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__a22o_1 _11124_ (.A1(\r1.regblock[16][19] ),
    .A2(_05860_),
    .B1(_05861_),
    .B2(_05863_),
    .X(_02640_));
 sky130_fd_sc_hd__clkbuf_1 _11125_ (.A(_05857_),
    .X(_01614_));
 sky130_fd_sc_hd__buf_1 _11126_ (.A(_05669_),
    .X(_05864_));
 sky130_fd_sc_hd__a22o_1 _11127_ (.A1(\r1.regblock[16][18] ),
    .A2(_05860_),
    .B1(_05864_),
    .B2(_05863_),
    .X(_02639_));
 sky130_fd_sc_hd__buf_2 _11128_ (.A(_05850_),
    .X(_05865_));
 sky130_fd_sc_hd__clkbuf_1 _11129_ (.A(_05865_),
    .X(_01613_));
 sky130_fd_sc_hd__buf_1 _11130_ (.A(_05673_),
    .X(_05866_));
 sky130_fd_sc_hd__a22o_1 _11131_ (.A1(\r1.regblock[16][17] ),
    .A2(_05860_),
    .B1(_05866_),
    .B2(_05863_),
    .X(_02638_));
 sky130_fd_sc_hd__clkbuf_1 _11132_ (.A(_05865_),
    .X(_01612_));
 sky130_fd_sc_hd__buf_1 _11133_ (.A(_05859_),
    .X(_05867_));
 sky130_fd_sc_hd__buf_1 _11134_ (.A(_05676_),
    .X(_05868_));
 sky130_fd_sc_hd__buf_1 _11135_ (.A(_05862_),
    .X(_05869_));
 sky130_fd_sc_hd__a22o_1 _11136_ (.A1(\r1.regblock[16][16] ),
    .A2(_05867_),
    .B1(_05868_),
    .B2(_05869_),
    .X(_02637_));
 sky130_fd_sc_hd__clkbuf_1 _11137_ (.A(_05865_),
    .X(_01611_));
 sky130_fd_sc_hd__buf_1 _11138_ (.A(_05679_),
    .X(_05870_));
 sky130_fd_sc_hd__a22o_1 _11139_ (.A1(\r1.regblock[16][15] ),
    .A2(_05867_),
    .B1(_05870_),
    .B2(_05869_),
    .X(_02636_));
 sky130_fd_sc_hd__clkbuf_2 _11140_ (.A(_05770_),
    .X(_05871_));
 sky130_fd_sc_hd__buf_2 _11141_ (.A(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__buf_1 _11142_ (.A(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__clkbuf_1 _11143_ (.A(_05873_),
    .X(_01610_));
 sky130_fd_sc_hd__buf_1 _11144_ (.A(_05682_),
    .X(_05874_));
 sky130_fd_sc_hd__a22o_1 _11145_ (.A1(\r1.regblock[16][14] ),
    .A2(_05867_),
    .B1(_05874_),
    .B2(_05869_),
    .X(_02635_));
 sky130_fd_sc_hd__clkbuf_1 _11146_ (.A(_05873_),
    .X(_01609_));
 sky130_fd_sc_hd__buf_1 _11147_ (.A(_05859_),
    .X(_05875_));
 sky130_fd_sc_hd__buf_1 _11148_ (.A(_05685_),
    .X(_05876_));
 sky130_fd_sc_hd__buf_1 _11149_ (.A(_05862_),
    .X(_05877_));
 sky130_fd_sc_hd__a22o_1 _11150_ (.A1(\r1.regblock[16][13] ),
    .A2(_05875_),
    .B1(_05876_),
    .B2(_05877_),
    .X(_02634_));
 sky130_fd_sc_hd__clkbuf_1 _11151_ (.A(_05873_),
    .X(_01608_));
 sky130_fd_sc_hd__buf_1 _11152_ (.A(_05688_),
    .X(_05878_));
 sky130_fd_sc_hd__a22o_1 _11153_ (.A1(\r1.regblock[16][12] ),
    .A2(_05875_),
    .B1(_05878_),
    .B2(_05877_),
    .X(_02633_));
 sky130_fd_sc_hd__buf_2 _11154_ (.A(_05872_),
    .X(_05879_));
 sky130_fd_sc_hd__clkbuf_1 _11155_ (.A(_05879_),
    .X(_01607_));
 sky130_fd_sc_hd__buf_1 _11156_ (.A(_05691_),
    .X(_05880_));
 sky130_fd_sc_hd__a22o_1 _11157_ (.A1(\r1.regblock[16][11] ),
    .A2(_05875_),
    .B1(_05880_),
    .B2(_05877_),
    .X(_02632_));
 sky130_fd_sc_hd__clkbuf_1 _11158_ (.A(_05879_),
    .X(_01606_));
 sky130_fd_sc_hd__buf_1 _11159_ (.A(_05836_),
    .X(_05881_));
 sky130_fd_sc_hd__buf_1 _11160_ (.A(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__buf_1 _11161_ (.A(_05695_),
    .X(_05883_));
 sky130_fd_sc_hd__buf_1 _11162_ (.A(_05840_),
    .X(_05884_));
 sky130_fd_sc_hd__buf_1 _11163_ (.A(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__a22o_1 _11164_ (.A1(\r1.regblock[16][10] ),
    .A2(_05882_),
    .B1(_05883_),
    .B2(_05885_),
    .X(_02631_));
 sky130_fd_sc_hd__clkbuf_1 _11165_ (.A(_05879_),
    .X(_01605_));
 sky130_fd_sc_hd__buf_1 _11166_ (.A(_05699_),
    .X(_05886_));
 sky130_fd_sc_hd__a22o_1 _11167_ (.A1(\r1.regblock[16][9] ),
    .A2(_05882_),
    .B1(_05886_),
    .B2(_05885_),
    .X(_02630_));
 sky130_fd_sc_hd__buf_1 _11168_ (.A(_05872_),
    .X(_05887_));
 sky130_fd_sc_hd__clkbuf_1 _11169_ (.A(_05887_),
    .X(_01604_));
 sky130_fd_sc_hd__buf_1 _11170_ (.A(_05703_),
    .X(_05888_));
 sky130_fd_sc_hd__a22o_1 _11171_ (.A1(\r1.regblock[16][8] ),
    .A2(_05882_),
    .B1(_05888_),
    .B2(_05885_),
    .X(_02629_));
 sky130_fd_sc_hd__clkbuf_1 _11172_ (.A(_05887_),
    .X(_01603_));
 sky130_fd_sc_hd__buf_1 _11173_ (.A(_05881_),
    .X(_05889_));
 sky130_fd_sc_hd__buf_1 _11174_ (.A(_05706_),
    .X(_05890_));
 sky130_fd_sc_hd__buf_1 _11175_ (.A(_05884_),
    .X(_05891_));
 sky130_fd_sc_hd__a22o_1 _11176_ (.A1(\r1.regblock[16][7] ),
    .A2(_05889_),
    .B1(_05890_),
    .B2(_05891_),
    .X(_02628_));
 sky130_fd_sc_hd__clkbuf_1 _11177_ (.A(_05887_),
    .X(_01602_));
 sky130_fd_sc_hd__buf_1 _11178_ (.A(_05709_),
    .X(_05892_));
 sky130_fd_sc_hd__a22o_1 _11179_ (.A1(\r1.regblock[16][6] ),
    .A2(_05889_),
    .B1(_05892_),
    .B2(_05891_),
    .X(_02627_));
 sky130_fd_sc_hd__clkbuf_2 _11180_ (.A(_05871_),
    .X(_05893_));
 sky130_fd_sc_hd__buf_1 _11181_ (.A(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__clkbuf_1 _11182_ (.A(_05894_),
    .X(_01601_));
 sky130_fd_sc_hd__buf_1 _11183_ (.A(_05712_),
    .X(_05895_));
 sky130_fd_sc_hd__a22o_1 _11184_ (.A1(\r1.regblock[16][5] ),
    .A2(_05889_),
    .B1(_05895_),
    .B2(_05891_),
    .X(_02626_));
 sky130_fd_sc_hd__clkbuf_1 _11185_ (.A(_05894_),
    .X(_01600_));
 sky130_fd_sc_hd__buf_1 _11186_ (.A(_05881_),
    .X(_05896_));
 sky130_fd_sc_hd__buf_1 _11187_ (.A(_05715_),
    .X(_05897_));
 sky130_fd_sc_hd__buf_1 _11188_ (.A(_05884_),
    .X(_05898_));
 sky130_fd_sc_hd__a22o_1 _11189_ (.A1(\r1.regblock[16][4] ),
    .A2(_05896_),
    .B1(_05897_),
    .B2(_05898_),
    .X(_02625_));
 sky130_fd_sc_hd__clkbuf_1 _11190_ (.A(_05894_),
    .X(_01599_));
 sky130_fd_sc_hd__buf_1 _11191_ (.A(_05718_),
    .X(_05899_));
 sky130_fd_sc_hd__a22o_1 _11192_ (.A1(\r1.regblock[16][3] ),
    .A2(_05896_),
    .B1(_05899_),
    .B2(_05898_),
    .X(_02624_));
 sky130_fd_sc_hd__buf_1 _11193_ (.A(_05893_),
    .X(_05900_));
 sky130_fd_sc_hd__clkbuf_1 _11194_ (.A(_05900_),
    .X(_01598_));
 sky130_fd_sc_hd__buf_1 _11195_ (.A(_05721_),
    .X(_05901_));
 sky130_fd_sc_hd__a22o_1 _11196_ (.A1(\r1.regblock[16][2] ),
    .A2(_05896_),
    .B1(_05901_),
    .B2(_05898_),
    .X(_02623_));
 sky130_fd_sc_hd__clkbuf_1 _11197_ (.A(_05900_),
    .X(_01597_));
 sky130_fd_sc_hd__buf_1 _11198_ (.A(_05723_),
    .X(_05902_));
 sky130_fd_sc_hd__a22o_1 _11199_ (.A1(\r1.regblock[16][1] ),
    .A2(_05827_),
    .B1(_05902_),
    .B2(_05831_),
    .X(_02622_));
 sky130_fd_sc_hd__clkbuf_1 _11200_ (.A(_05900_),
    .X(_01596_));
 sky130_fd_sc_hd__buf_1 _11201_ (.A(_05725_),
    .X(_05903_));
 sky130_fd_sc_hd__a22o_1 _11202_ (.A1(\r1.regblock[16][0] ),
    .A2(_05827_),
    .B1(_05903_),
    .B2(_05831_),
    .X(_02621_));
 sky130_fd_sc_hd__buf_1 _11203_ (.A(_05893_),
    .X(_05904_));
 sky130_fd_sc_hd__clkbuf_1 _11204_ (.A(_05904_),
    .X(_01595_));
 sky130_fd_sc_hd__or2_2 _11205_ (.A(_05825_),
    .B(_04640_),
    .X(_05905_));
 sky130_fd_sc_hd__buf_1 _11206_ (.A(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__buf_1 _11207_ (.A(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__inv_2 _11208_ (.A(_05905_),
    .Y(_05908_));
 sky130_fd_sc_hd__buf_1 _11209_ (.A(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__buf_1 _11210_ (.A(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__a22o_1 _11211_ (.A1(\r1.regblock[17][31] ),
    .A2(_05907_),
    .B1(_05829_),
    .B2(_05910_),
    .X(_02620_));
 sky130_fd_sc_hd__clkbuf_1 _11212_ (.A(_05904_),
    .X(_01594_));
 sky130_fd_sc_hd__a22o_1 _11213_ (.A1(\r1.regblock[17][30] ),
    .A2(_05907_),
    .B1(_05833_),
    .B2(_05910_),
    .X(_02619_));
 sky130_fd_sc_hd__clkbuf_1 _11214_ (.A(_05904_),
    .X(_01593_));
 sky130_fd_sc_hd__a22o_1 _11215_ (.A1(\r1.regblock[17][29] ),
    .A2(_05907_),
    .B1(_05835_),
    .B2(_05910_),
    .X(_02618_));
 sky130_fd_sc_hd__buf_2 _11216_ (.A(_05871_),
    .X(_05911_));
 sky130_fd_sc_hd__buf_1 _11217_ (.A(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__clkbuf_1 _11218_ (.A(_05912_),
    .X(_01592_));
 sky130_fd_sc_hd__buf_2 _11219_ (.A(_05905_),
    .X(_05913_));
 sky130_fd_sc_hd__buf_2 _11220_ (.A(_05913_),
    .X(_05914_));
 sky130_fd_sc_hd__buf_1 _11221_ (.A(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__buf_2 _11222_ (.A(_05908_),
    .X(_05916_));
 sky130_fd_sc_hd__buf_2 _11223_ (.A(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__buf_1 _11224_ (.A(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__a22o_1 _11225_ (.A1(\r1.regblock[17][28] ),
    .A2(_05915_),
    .B1(_05839_),
    .B2(_05918_),
    .X(_02617_));
 sky130_fd_sc_hd__clkbuf_1 _11226_ (.A(_05912_),
    .X(_01591_));
 sky130_fd_sc_hd__a22o_1 _11227_ (.A1(\r1.regblock[17][27] ),
    .A2(_05915_),
    .B1(_05843_),
    .B2(_05918_),
    .X(_02616_));
 sky130_fd_sc_hd__clkbuf_1 _11228_ (.A(_05912_),
    .X(_01590_));
 sky130_fd_sc_hd__a22o_1 _11229_ (.A1(\r1.regblock[17][26] ),
    .A2(_05915_),
    .B1(_05845_),
    .B2(_05918_),
    .X(_02615_));
 sky130_fd_sc_hd__buf_1 _11230_ (.A(_05911_),
    .X(_05919_));
 sky130_fd_sc_hd__clkbuf_1 _11231_ (.A(_05919_),
    .X(_01589_));
 sky130_fd_sc_hd__buf_1 _11232_ (.A(_05914_),
    .X(_05920_));
 sky130_fd_sc_hd__buf_1 _11233_ (.A(_05917_),
    .X(_05921_));
 sky130_fd_sc_hd__a22o_1 _11234_ (.A1(\r1.regblock[17][25] ),
    .A2(_05920_),
    .B1(_05847_),
    .B2(_05921_),
    .X(_02614_));
 sky130_fd_sc_hd__clkbuf_1 _11235_ (.A(_05919_),
    .X(_01588_));
 sky130_fd_sc_hd__a22o_1 _11236_ (.A1(\r1.regblock[17][24] ),
    .A2(_05920_),
    .B1(_05849_),
    .B2(_05921_),
    .X(_02613_));
 sky130_fd_sc_hd__clkbuf_1 _11237_ (.A(_05919_),
    .X(_01587_));
 sky130_fd_sc_hd__a22o_1 _11238_ (.A1(\r1.regblock[17][23] ),
    .A2(_05920_),
    .B1(_05852_),
    .B2(_05921_),
    .X(_02612_));
 sky130_fd_sc_hd__buf_1 _11239_ (.A(_05911_),
    .X(_05922_));
 sky130_fd_sc_hd__clkbuf_1 _11240_ (.A(_05922_),
    .X(_01586_));
 sky130_fd_sc_hd__buf_1 _11241_ (.A(_05914_),
    .X(_05923_));
 sky130_fd_sc_hd__buf_1 _11242_ (.A(_05917_),
    .X(_05924_));
 sky130_fd_sc_hd__a22o_1 _11243_ (.A1(\r1.regblock[17][22] ),
    .A2(_05923_),
    .B1(_05854_),
    .B2(_05924_),
    .X(_02611_));
 sky130_fd_sc_hd__clkbuf_1 _11244_ (.A(_05922_),
    .X(_01585_));
 sky130_fd_sc_hd__a22o_1 _11245_ (.A1(\r1.regblock[17][21] ),
    .A2(_05923_),
    .B1(_05856_),
    .B2(_05924_),
    .X(_02610_));
 sky130_fd_sc_hd__clkbuf_1 _11246_ (.A(_05922_),
    .X(_01584_));
 sky130_fd_sc_hd__a22o_1 _11247_ (.A1(\r1.regblock[17][20] ),
    .A2(_05923_),
    .B1(_05858_),
    .B2(_05924_),
    .X(_02609_));
 sky130_fd_sc_hd__clkbuf_1 _11248_ (.A(_03907_),
    .X(_05925_));
 sky130_fd_sc_hd__buf_1 _11249_ (.A(_05925_),
    .X(_05926_));
 sky130_fd_sc_hd__buf_2 _11250_ (.A(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__buf_1 _11251_ (.A(_05927_),
    .X(_05928_));
 sky130_fd_sc_hd__clkbuf_1 _11252_ (.A(_05928_),
    .X(_01583_));
 sky130_fd_sc_hd__buf_2 _11253_ (.A(_05913_),
    .X(_05929_));
 sky130_fd_sc_hd__buf_1 _11254_ (.A(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__buf_2 _11255_ (.A(_05916_),
    .X(_05931_));
 sky130_fd_sc_hd__buf_1 _11256_ (.A(_05931_),
    .X(_05932_));
 sky130_fd_sc_hd__a22o_1 _11257_ (.A1(\r1.regblock[17][19] ),
    .A2(_05930_),
    .B1(_05861_),
    .B2(_05932_),
    .X(_02608_));
 sky130_fd_sc_hd__clkbuf_1 _11258_ (.A(_05928_),
    .X(_01582_));
 sky130_fd_sc_hd__a22o_1 _11259_ (.A1(\r1.regblock[17][18] ),
    .A2(_05930_),
    .B1(_05864_),
    .B2(_05932_),
    .X(_02607_));
 sky130_fd_sc_hd__clkbuf_1 _11260_ (.A(_05928_),
    .X(_01581_));
 sky130_fd_sc_hd__a22o_1 _11261_ (.A1(\r1.regblock[17][17] ),
    .A2(_05930_),
    .B1(_05866_),
    .B2(_05932_),
    .X(_02606_));
 sky130_fd_sc_hd__buf_1 _11262_ (.A(_05927_),
    .X(_05933_));
 sky130_fd_sc_hd__clkbuf_1 _11263_ (.A(_05933_),
    .X(_01580_));
 sky130_fd_sc_hd__buf_1 _11264_ (.A(_05929_),
    .X(_05934_));
 sky130_fd_sc_hd__buf_1 _11265_ (.A(_05931_),
    .X(_05935_));
 sky130_fd_sc_hd__a22o_1 _11266_ (.A1(\r1.regblock[17][16] ),
    .A2(_05934_),
    .B1(_05868_),
    .B2(_05935_),
    .X(_02605_));
 sky130_fd_sc_hd__clkbuf_1 _11267_ (.A(_05933_),
    .X(_01579_));
 sky130_fd_sc_hd__a22o_1 _11268_ (.A1(\r1.regblock[17][15] ),
    .A2(_05934_),
    .B1(_05870_),
    .B2(_05935_),
    .X(_02604_));
 sky130_fd_sc_hd__clkbuf_1 _11269_ (.A(_05933_),
    .X(_01578_));
 sky130_fd_sc_hd__a22o_1 _11270_ (.A1(\r1.regblock[17][14] ),
    .A2(_05934_),
    .B1(_05874_),
    .B2(_05935_),
    .X(_02603_));
 sky130_fd_sc_hd__buf_1 _11271_ (.A(_05927_),
    .X(_05936_));
 sky130_fd_sc_hd__clkbuf_1 _11272_ (.A(_05936_),
    .X(_01577_));
 sky130_fd_sc_hd__buf_1 _11273_ (.A(_05929_),
    .X(_05937_));
 sky130_fd_sc_hd__buf_1 _11274_ (.A(_05931_),
    .X(_05938_));
 sky130_fd_sc_hd__a22o_1 _11275_ (.A1(\r1.regblock[17][13] ),
    .A2(_05937_),
    .B1(_05876_),
    .B2(_05938_),
    .X(_02602_));
 sky130_fd_sc_hd__clkbuf_1 _11276_ (.A(_05936_),
    .X(_01576_));
 sky130_fd_sc_hd__a22o_1 _11277_ (.A1(\r1.regblock[17][12] ),
    .A2(_05937_),
    .B1(_05878_),
    .B2(_05938_),
    .X(_02601_));
 sky130_fd_sc_hd__clkbuf_1 _11278_ (.A(_05936_),
    .X(_01575_));
 sky130_fd_sc_hd__a22o_1 _11279_ (.A1(\r1.regblock[17][11] ),
    .A2(_05937_),
    .B1(_05880_),
    .B2(_05938_),
    .X(_02600_));
 sky130_fd_sc_hd__clkbuf_2 _11280_ (.A(_05926_),
    .X(_05939_));
 sky130_fd_sc_hd__buf_1 _11281_ (.A(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__clkbuf_1 _11282_ (.A(_05940_),
    .X(_01574_));
 sky130_fd_sc_hd__clkbuf_2 _11283_ (.A(_05913_),
    .X(_05941_));
 sky130_fd_sc_hd__buf_1 _11284_ (.A(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__clkbuf_2 _11285_ (.A(_05916_),
    .X(_05943_));
 sky130_fd_sc_hd__buf_1 _11286_ (.A(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__a22o_1 _11287_ (.A1(\r1.regblock[17][10] ),
    .A2(_05942_),
    .B1(_05883_),
    .B2(_05944_),
    .X(_02599_));
 sky130_fd_sc_hd__clkbuf_1 _11288_ (.A(_05940_),
    .X(_01573_));
 sky130_fd_sc_hd__a22o_1 _11289_ (.A1(\r1.regblock[17][9] ),
    .A2(_05942_),
    .B1(_05886_),
    .B2(_05944_),
    .X(_02598_));
 sky130_fd_sc_hd__clkbuf_1 _11290_ (.A(_05940_),
    .X(_01572_));
 sky130_fd_sc_hd__a22o_1 _11291_ (.A1(\r1.regblock[17][8] ),
    .A2(_05942_),
    .B1(_05888_),
    .B2(_05944_),
    .X(_02597_));
 sky130_fd_sc_hd__buf_1 _11292_ (.A(_05939_),
    .X(_05945_));
 sky130_fd_sc_hd__clkbuf_1 _11293_ (.A(_05945_),
    .X(_01571_));
 sky130_fd_sc_hd__buf_1 _11294_ (.A(_05941_),
    .X(_05946_));
 sky130_fd_sc_hd__buf_1 _11295_ (.A(_05943_),
    .X(_05947_));
 sky130_fd_sc_hd__a22o_1 _11296_ (.A1(\r1.regblock[17][7] ),
    .A2(_05946_),
    .B1(_05890_),
    .B2(_05947_),
    .X(_02596_));
 sky130_fd_sc_hd__clkbuf_1 _11297_ (.A(_05945_),
    .X(_01570_));
 sky130_fd_sc_hd__a22o_1 _11298_ (.A1(\r1.regblock[17][6] ),
    .A2(_05946_),
    .B1(_05892_),
    .B2(_05947_),
    .X(_02595_));
 sky130_fd_sc_hd__clkbuf_1 _11299_ (.A(_05945_),
    .X(_01569_));
 sky130_fd_sc_hd__a22o_1 _11300_ (.A1(\r1.regblock[17][5] ),
    .A2(_05946_),
    .B1(_05895_),
    .B2(_05947_),
    .X(_02594_));
 sky130_fd_sc_hd__buf_1 _11301_ (.A(_05939_),
    .X(_05948_));
 sky130_fd_sc_hd__clkbuf_1 _11302_ (.A(_05948_),
    .X(_01568_));
 sky130_fd_sc_hd__buf_1 _11303_ (.A(_05941_),
    .X(_05949_));
 sky130_fd_sc_hd__buf_1 _11304_ (.A(_05943_),
    .X(_05950_));
 sky130_fd_sc_hd__a22o_1 _11305_ (.A1(\r1.regblock[17][4] ),
    .A2(_05949_),
    .B1(_05897_),
    .B2(_05950_),
    .X(_02593_));
 sky130_fd_sc_hd__clkbuf_1 _11306_ (.A(_05948_),
    .X(_01567_));
 sky130_fd_sc_hd__a22o_1 _11307_ (.A1(\r1.regblock[17][3] ),
    .A2(_05949_),
    .B1(_05899_),
    .B2(_05950_),
    .X(_02592_));
 sky130_fd_sc_hd__clkbuf_1 _11308_ (.A(_05948_),
    .X(_01566_));
 sky130_fd_sc_hd__a22o_1 _11309_ (.A1(\r1.regblock[17][2] ),
    .A2(_05949_),
    .B1(_05901_),
    .B2(_05950_),
    .X(_02591_));
 sky130_fd_sc_hd__buf_2 _11310_ (.A(_05926_),
    .X(_05951_));
 sky130_fd_sc_hd__buf_1 _11311_ (.A(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__clkbuf_1 _11312_ (.A(_05952_),
    .X(_01565_));
 sky130_fd_sc_hd__a22o_1 _11313_ (.A1(\r1.regblock[17][1] ),
    .A2(_05906_),
    .B1(_05902_),
    .B2(_05909_),
    .X(_02590_));
 sky130_fd_sc_hd__clkbuf_1 _11314_ (.A(_05952_),
    .X(_01564_));
 sky130_fd_sc_hd__a22o_1 _11315_ (.A1(\r1.regblock[17][0] ),
    .A2(_05906_),
    .B1(_05903_),
    .B2(_05909_),
    .X(_02589_));
 sky130_fd_sc_hd__clkbuf_1 _11316_ (.A(_05952_),
    .X(_01563_));
 sky130_fd_sc_hd__or2_2 _11317_ (.A(_05825_),
    .B(_05053_),
    .X(_05953_));
 sky130_fd_sc_hd__buf_1 _11318_ (.A(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__buf_1 _11319_ (.A(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__inv_2 _11320_ (.A(_05953_),
    .Y(_05956_));
 sky130_fd_sc_hd__buf_1 _11321_ (.A(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__buf_1 _11322_ (.A(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__a22o_1 _11323_ (.A1(\r1.regblock[18][31] ),
    .A2(_05955_),
    .B1(_05829_),
    .B2(_05958_),
    .X(_02588_));
 sky130_fd_sc_hd__buf_1 _11324_ (.A(_05951_),
    .X(_05959_));
 sky130_fd_sc_hd__clkbuf_1 _11325_ (.A(_05959_),
    .X(_01562_));
 sky130_fd_sc_hd__a22o_1 _11326_ (.A1(\r1.regblock[18][30] ),
    .A2(_05955_),
    .B1(_05833_),
    .B2(_05958_),
    .X(_02587_));
 sky130_fd_sc_hd__clkbuf_1 _11327_ (.A(_05959_),
    .X(_01561_));
 sky130_fd_sc_hd__a22o_1 _11328_ (.A1(\r1.regblock[18][29] ),
    .A2(_05955_),
    .B1(_05835_),
    .B2(_05958_),
    .X(_02586_));
 sky130_fd_sc_hd__clkbuf_1 _11329_ (.A(_05959_),
    .X(_01560_));
 sky130_fd_sc_hd__clkbuf_2 _11330_ (.A(_05953_),
    .X(_05960_));
 sky130_fd_sc_hd__buf_2 _11331_ (.A(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__buf_1 _11332_ (.A(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__buf_2 _11333_ (.A(_05956_),
    .X(_05963_));
 sky130_fd_sc_hd__buf_2 _11334_ (.A(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__buf_1 _11335_ (.A(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__a22o_1 _11336_ (.A1(\r1.regblock[18][28] ),
    .A2(_05962_),
    .B1(_05839_),
    .B2(_05965_),
    .X(_02585_));
 sky130_fd_sc_hd__buf_1 _11337_ (.A(_05951_),
    .X(_05966_));
 sky130_fd_sc_hd__clkbuf_1 _11338_ (.A(_05966_),
    .X(_01559_));
 sky130_fd_sc_hd__a22o_1 _11339_ (.A1(\r1.regblock[18][27] ),
    .A2(_05962_),
    .B1(_05843_),
    .B2(_05965_),
    .X(_02584_));
 sky130_fd_sc_hd__clkbuf_1 _11340_ (.A(_05966_),
    .X(_01558_));
 sky130_fd_sc_hd__a22o_1 _11341_ (.A1(\r1.regblock[18][26] ),
    .A2(_05962_),
    .B1(_05845_),
    .B2(_05965_),
    .X(_02583_));
 sky130_fd_sc_hd__clkbuf_1 _11342_ (.A(_05966_),
    .X(_01557_));
 sky130_fd_sc_hd__buf_1 _11343_ (.A(_05961_),
    .X(_05967_));
 sky130_fd_sc_hd__buf_1 _11344_ (.A(_05964_),
    .X(_05968_));
 sky130_fd_sc_hd__a22o_1 _11345_ (.A1(\r1.regblock[18][25] ),
    .A2(_05967_),
    .B1(_05847_),
    .B2(_05968_),
    .X(_02582_));
 sky130_fd_sc_hd__buf_1 _11346_ (.A(_05925_),
    .X(_05969_));
 sky130_fd_sc_hd__clkbuf_2 _11347_ (.A(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__buf_2 _11348_ (.A(_05970_),
    .X(_05971_));
 sky130_fd_sc_hd__clkbuf_1 _11349_ (.A(_05971_),
    .X(_01556_));
 sky130_fd_sc_hd__a22o_1 _11350_ (.A1(\r1.regblock[18][24] ),
    .A2(_05967_),
    .B1(_05849_),
    .B2(_05968_),
    .X(_02581_));
 sky130_fd_sc_hd__clkbuf_1 _11351_ (.A(_05971_),
    .X(_01555_));
 sky130_fd_sc_hd__a22o_1 _11352_ (.A1(\r1.regblock[18][23] ),
    .A2(_05967_),
    .B1(_05852_),
    .B2(_05968_),
    .X(_02580_));
 sky130_fd_sc_hd__clkbuf_1 _11353_ (.A(_05971_),
    .X(_01554_));
 sky130_fd_sc_hd__buf_1 _11354_ (.A(_05961_),
    .X(_05972_));
 sky130_fd_sc_hd__buf_1 _11355_ (.A(_05964_),
    .X(_05973_));
 sky130_fd_sc_hd__a22o_1 _11356_ (.A1(\r1.regblock[18][22] ),
    .A2(_05972_),
    .B1(_05854_),
    .B2(_05973_),
    .X(_02579_));
 sky130_fd_sc_hd__buf_2 _11357_ (.A(_05970_),
    .X(_05974_));
 sky130_fd_sc_hd__clkbuf_1 _11358_ (.A(_05974_),
    .X(_01553_));
 sky130_fd_sc_hd__a22o_1 _11359_ (.A1(\r1.regblock[18][21] ),
    .A2(_05972_),
    .B1(_05856_),
    .B2(_05973_),
    .X(_02578_));
 sky130_fd_sc_hd__clkbuf_1 _11360_ (.A(_05974_),
    .X(_01552_));
 sky130_fd_sc_hd__a22o_1 _11361_ (.A1(\r1.regblock[18][20] ),
    .A2(_05972_),
    .B1(_05858_),
    .B2(_05973_),
    .X(_02577_));
 sky130_fd_sc_hd__clkbuf_1 _11362_ (.A(_05974_),
    .X(_01551_));
 sky130_fd_sc_hd__buf_2 _11363_ (.A(_05960_),
    .X(_05975_));
 sky130_fd_sc_hd__buf_1 _11364_ (.A(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__buf_2 _11365_ (.A(_05963_),
    .X(_05977_));
 sky130_fd_sc_hd__buf_1 _11366_ (.A(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__a22o_1 _11367_ (.A1(\r1.regblock[18][19] ),
    .A2(_05976_),
    .B1(_05861_),
    .B2(_05978_),
    .X(_02576_));
 sky130_fd_sc_hd__buf_2 _11368_ (.A(_05970_),
    .X(_05979_));
 sky130_fd_sc_hd__clkbuf_1 _11369_ (.A(_05979_),
    .X(_01550_));
 sky130_fd_sc_hd__a22o_1 _11370_ (.A1(\r1.regblock[18][18] ),
    .A2(_05976_),
    .B1(_05864_),
    .B2(_05978_),
    .X(_02575_));
 sky130_fd_sc_hd__clkbuf_1 _11371_ (.A(_05979_),
    .X(_01549_));
 sky130_fd_sc_hd__a22o_1 _11372_ (.A1(\r1.regblock[18][17] ),
    .A2(_05976_),
    .B1(_05866_),
    .B2(_05978_),
    .X(_02574_));
 sky130_fd_sc_hd__clkbuf_1 _11373_ (.A(_05979_),
    .X(_01548_));
 sky130_fd_sc_hd__buf_1 _11374_ (.A(_05975_),
    .X(_05980_));
 sky130_fd_sc_hd__buf_1 _11375_ (.A(_05977_),
    .X(_05981_));
 sky130_fd_sc_hd__a22o_1 _11376_ (.A1(\r1.regblock[18][16] ),
    .A2(_05980_),
    .B1(_05868_),
    .B2(_05981_),
    .X(_02573_));
 sky130_fd_sc_hd__clkbuf_4 _11377_ (.A(_05969_),
    .X(_05982_));
 sky130_fd_sc_hd__buf_1 _11378_ (.A(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__clkbuf_1 _11379_ (.A(_05983_),
    .X(_01547_));
 sky130_fd_sc_hd__a22o_1 _11380_ (.A1(\r1.regblock[18][15] ),
    .A2(_05980_),
    .B1(_05870_),
    .B2(_05981_),
    .X(_02572_));
 sky130_fd_sc_hd__clkbuf_1 _11381_ (.A(_05983_),
    .X(_01546_));
 sky130_fd_sc_hd__a22o_1 _11382_ (.A1(\r1.regblock[18][14] ),
    .A2(_05980_),
    .B1(_05874_),
    .B2(_05981_),
    .X(_02571_));
 sky130_fd_sc_hd__clkbuf_1 _11383_ (.A(_05983_),
    .X(_01545_));
 sky130_fd_sc_hd__buf_1 _11384_ (.A(_05975_),
    .X(_05984_));
 sky130_fd_sc_hd__buf_1 _11385_ (.A(_05977_),
    .X(_05985_));
 sky130_fd_sc_hd__a22o_1 _11386_ (.A1(\r1.regblock[18][13] ),
    .A2(_05984_),
    .B1(_05876_),
    .B2(_05985_),
    .X(_02570_));
 sky130_fd_sc_hd__buf_2 _11387_ (.A(_05982_),
    .X(_05986_));
 sky130_fd_sc_hd__clkbuf_1 _11388_ (.A(_05986_),
    .X(_01544_));
 sky130_fd_sc_hd__a22o_1 _11389_ (.A1(\r1.regblock[18][12] ),
    .A2(_05984_),
    .B1(_05878_),
    .B2(_05985_),
    .X(_02569_));
 sky130_fd_sc_hd__clkbuf_1 _11390_ (.A(_05986_),
    .X(_01543_));
 sky130_fd_sc_hd__a22o_1 _11391_ (.A1(\r1.regblock[18][11] ),
    .A2(_05984_),
    .B1(_05880_),
    .B2(_05985_),
    .X(_02568_));
 sky130_fd_sc_hd__clkbuf_1 _11392_ (.A(_05986_),
    .X(_01542_));
 sky130_fd_sc_hd__clkbuf_2 _11393_ (.A(_05960_),
    .X(_05987_));
 sky130_fd_sc_hd__buf_1 _11394_ (.A(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__clkbuf_2 _11395_ (.A(_05963_),
    .X(_05989_));
 sky130_fd_sc_hd__buf_1 _11396_ (.A(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__a22o_1 _11397_ (.A1(\r1.regblock[18][10] ),
    .A2(_05988_),
    .B1(_05883_),
    .B2(_05990_),
    .X(_02567_));
 sky130_fd_sc_hd__buf_1 _11398_ (.A(_05982_),
    .X(_05991_));
 sky130_fd_sc_hd__clkbuf_1 _11399_ (.A(_05991_),
    .X(_01541_));
 sky130_fd_sc_hd__a22o_1 _11400_ (.A1(\r1.regblock[18][9] ),
    .A2(_05988_),
    .B1(_05886_),
    .B2(_05990_),
    .X(_02566_));
 sky130_fd_sc_hd__clkbuf_1 _11401_ (.A(_05991_),
    .X(_01540_));
 sky130_fd_sc_hd__a22o_1 _11402_ (.A1(\r1.regblock[18][8] ),
    .A2(_05988_),
    .B1(_05888_),
    .B2(_05990_),
    .X(_02565_));
 sky130_fd_sc_hd__clkbuf_1 _11403_ (.A(_05991_),
    .X(_01539_));
 sky130_fd_sc_hd__buf_1 _11404_ (.A(_05987_),
    .X(_05992_));
 sky130_fd_sc_hd__buf_1 _11405_ (.A(_05989_),
    .X(_05993_));
 sky130_fd_sc_hd__a22o_1 _11406_ (.A1(\r1.regblock[18][7] ),
    .A2(_05992_),
    .B1(_05890_),
    .B2(_05993_),
    .X(_02564_));
 sky130_fd_sc_hd__buf_1 _11407_ (.A(_05969_),
    .X(_05994_));
 sky130_fd_sc_hd__buf_1 _11408_ (.A(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__clkbuf_1 _11409_ (.A(_05995_),
    .X(_01538_));
 sky130_fd_sc_hd__a22o_1 _11410_ (.A1(\r1.regblock[18][6] ),
    .A2(_05992_),
    .B1(_05892_),
    .B2(_05993_),
    .X(_02563_));
 sky130_fd_sc_hd__clkbuf_1 _11411_ (.A(_05995_),
    .X(_01537_));
 sky130_fd_sc_hd__a22o_1 _11412_ (.A1(\r1.regblock[18][5] ),
    .A2(_05992_),
    .B1(_05895_),
    .B2(_05993_),
    .X(_02562_));
 sky130_fd_sc_hd__clkbuf_1 _11413_ (.A(_05995_),
    .X(_01536_));
 sky130_fd_sc_hd__buf_1 _11414_ (.A(_05987_),
    .X(_05996_));
 sky130_fd_sc_hd__buf_1 _11415_ (.A(_05989_),
    .X(_05997_));
 sky130_fd_sc_hd__a22o_1 _11416_ (.A1(\r1.regblock[18][4] ),
    .A2(_05996_),
    .B1(_05897_),
    .B2(_05997_),
    .X(_02561_));
 sky130_fd_sc_hd__buf_1 _11417_ (.A(_05994_),
    .X(_05998_));
 sky130_fd_sc_hd__clkbuf_1 _11418_ (.A(_05998_),
    .X(_01535_));
 sky130_fd_sc_hd__a22o_1 _11419_ (.A1(\r1.regblock[18][3] ),
    .A2(_05996_),
    .B1(_05899_),
    .B2(_05997_),
    .X(_02560_));
 sky130_fd_sc_hd__clkbuf_1 _11420_ (.A(_05998_),
    .X(_01534_));
 sky130_fd_sc_hd__a22o_1 _11421_ (.A1(\r1.regblock[18][2] ),
    .A2(_05996_),
    .B1(_05901_),
    .B2(_05997_),
    .X(_02559_));
 sky130_fd_sc_hd__buf_1 _11422_ (.A(_05998_),
    .X(_01533_));
 sky130_fd_sc_hd__a22o_1 _11423_ (.A1(\r1.regblock[18][1] ),
    .A2(_05954_),
    .B1(_05902_),
    .B2(_05957_),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_2 _11424_ (.A(_05994_),
    .X(_05999_));
 sky130_fd_sc_hd__clkbuf_1 _11425_ (.A(_05999_),
    .X(_01532_));
 sky130_fd_sc_hd__a22o_1 _11426_ (.A1(\r1.regblock[18][0] ),
    .A2(_05954_),
    .B1(_05903_),
    .B2(_05957_),
    .X(_02557_));
 sky130_fd_sc_hd__clkbuf_1 _11427_ (.A(_05999_),
    .X(_01531_));
 sky130_fd_sc_hd__or2_2 _11428_ (.A(_04216_),
    .B(_04640_),
    .X(_06000_));
 sky130_fd_sc_hd__buf_1 _11429_ (.A(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__buf_1 _11430_ (.A(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__buf_1 _11431_ (.A(_05620_),
    .X(_06003_));
 sky130_fd_sc_hd__inv_2 _11432_ (.A(_06000_),
    .Y(_06004_));
 sky130_fd_sc_hd__buf_1 _11433_ (.A(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__buf_1 _11434_ (.A(_06005_),
    .X(_06006_));
 sky130_fd_sc_hd__a22o_1 _11435_ (.A1(\r1.regblock[1][31] ),
    .A2(_06002_),
    .B1(_06003_),
    .B2(_06006_),
    .X(_02556_));
 sky130_fd_sc_hd__clkbuf_1 _11436_ (.A(_05999_),
    .X(_01530_));
 sky130_fd_sc_hd__buf_1 _11437_ (.A(_05625_),
    .X(_06007_));
 sky130_fd_sc_hd__a22o_1 _11438_ (.A1(\r1.regblock[1][30] ),
    .A2(_06002_),
    .B1(_06007_),
    .B2(_06006_),
    .X(_02555_));
 sky130_fd_sc_hd__buf_2 _11439_ (.A(_05925_),
    .X(_06008_));
 sky130_fd_sc_hd__clkbuf_2 _11440_ (.A(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__buf_1 _11441_ (.A(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__buf_1 _11442_ (.A(_06010_),
    .X(_01529_));
 sky130_fd_sc_hd__buf_1 _11443_ (.A(_05628_),
    .X(_06011_));
 sky130_fd_sc_hd__a22o_1 _11444_ (.A1(\r1.regblock[1][29] ),
    .A2(_06002_),
    .B1(_06011_),
    .B2(_06006_),
    .X(_02554_));
 sky130_fd_sc_hd__clkbuf_1 _11445_ (.A(_06010_),
    .X(_01528_));
 sky130_fd_sc_hd__clkbuf_4 _11446_ (.A(_06000_),
    .X(_06012_));
 sky130_fd_sc_hd__clkbuf_2 _11447_ (.A(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__buf_1 _11448_ (.A(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__clkbuf_2 _11449_ (.A(_05633_),
    .X(_06015_));
 sky130_fd_sc_hd__clkbuf_4 _11450_ (.A(_06004_),
    .X(_06016_));
 sky130_fd_sc_hd__clkbuf_2 _11451_ (.A(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__buf_1 _11452_ (.A(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__a22o_1 _11453_ (.A1(\r1.regblock[1][28] ),
    .A2(_06014_),
    .B1(_06015_),
    .B2(_06018_),
    .X(_02553_));
 sky130_fd_sc_hd__clkbuf_1 _11454_ (.A(_06010_),
    .X(_01527_));
 sky130_fd_sc_hd__clkbuf_2 _11455_ (.A(_05638_),
    .X(_06019_));
 sky130_fd_sc_hd__a22o_1 _11456_ (.A1(\r1.regblock[1][27] ),
    .A2(_06014_),
    .B1(_06019_),
    .B2(_06018_),
    .X(_02552_));
 sky130_fd_sc_hd__buf_1 _11457_ (.A(_06009_),
    .X(_06020_));
 sky130_fd_sc_hd__clkbuf_1 _11458_ (.A(_06020_),
    .X(_01526_));
 sky130_fd_sc_hd__clkbuf_2 _11459_ (.A(_05643_),
    .X(_06021_));
 sky130_fd_sc_hd__a22o_1 _11460_ (.A1(\r1.regblock[1][26] ),
    .A2(_06014_),
    .B1(_06021_),
    .B2(_06018_),
    .X(_02551_));
 sky130_fd_sc_hd__clkbuf_1 _11461_ (.A(_06020_),
    .X(_01525_));
 sky130_fd_sc_hd__buf_1 _11462_ (.A(_06013_),
    .X(_06022_));
 sky130_fd_sc_hd__buf_1 _11463_ (.A(_05646_),
    .X(_06023_));
 sky130_fd_sc_hd__buf_1 _11464_ (.A(_06017_),
    .X(_06024_));
 sky130_fd_sc_hd__a22o_1 _11465_ (.A1(\r1.regblock[1][25] ),
    .A2(_06022_),
    .B1(_06023_),
    .B2(_06024_),
    .X(_02550_));
 sky130_fd_sc_hd__clkbuf_1 _11466_ (.A(_06020_),
    .X(_01524_));
 sky130_fd_sc_hd__buf_1 _11467_ (.A(_05649_),
    .X(_06025_));
 sky130_fd_sc_hd__a22o_1 _11468_ (.A1(\r1.regblock[1][24] ),
    .A2(_06022_),
    .B1(_06025_),
    .B2(_06024_),
    .X(_02549_));
 sky130_fd_sc_hd__buf_1 _11469_ (.A(_06009_),
    .X(_06026_));
 sky130_fd_sc_hd__clkbuf_1 _11470_ (.A(_06026_),
    .X(_01523_));
 sky130_fd_sc_hd__buf_1 _11471_ (.A(_05652_),
    .X(_06027_));
 sky130_fd_sc_hd__a22o_1 _11472_ (.A1(\r1.regblock[1][23] ),
    .A2(_06022_),
    .B1(_06027_),
    .B2(_06024_),
    .X(_02548_));
 sky130_fd_sc_hd__clkbuf_1 _11473_ (.A(_06026_),
    .X(_01522_));
 sky130_fd_sc_hd__buf_1 _11474_ (.A(_06013_),
    .X(_06028_));
 sky130_fd_sc_hd__buf_1 _11475_ (.A(_05655_),
    .X(_06029_));
 sky130_fd_sc_hd__buf_1 _11476_ (.A(_06017_),
    .X(_06030_));
 sky130_fd_sc_hd__a22o_1 _11477_ (.A1(\r1.regblock[1][22] ),
    .A2(_06028_),
    .B1(_06029_),
    .B2(_06030_),
    .X(_02547_));
 sky130_fd_sc_hd__clkbuf_1 _11478_ (.A(_06026_),
    .X(_01521_));
 sky130_fd_sc_hd__buf_1 _11479_ (.A(_05658_),
    .X(_06031_));
 sky130_fd_sc_hd__a22o_1 _11480_ (.A1(\r1.regblock[1][21] ),
    .A2(_06028_),
    .B1(_06031_),
    .B2(_06030_),
    .X(_02546_));
 sky130_fd_sc_hd__clkbuf_2 _11481_ (.A(_06008_),
    .X(_06032_));
 sky130_fd_sc_hd__buf_1 _11482_ (.A(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__clkbuf_2 _11483_ (.A(_06033_),
    .X(_01520_));
 sky130_fd_sc_hd__buf_1 _11484_ (.A(_05661_),
    .X(_06034_));
 sky130_fd_sc_hd__a22o_1 _11485_ (.A1(\r1.regblock[1][20] ),
    .A2(_06028_),
    .B1(_06034_),
    .B2(_06030_),
    .X(_02545_));
 sky130_fd_sc_hd__clkbuf_1 _11486_ (.A(_06033_),
    .X(_01519_));
 sky130_fd_sc_hd__clkbuf_2 _11487_ (.A(_06012_),
    .X(_06035_));
 sky130_fd_sc_hd__buf_1 _11488_ (.A(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__buf_1 _11489_ (.A(_05665_),
    .X(_06037_));
 sky130_fd_sc_hd__clkbuf_2 _11490_ (.A(_06016_),
    .X(_06038_));
 sky130_fd_sc_hd__buf_1 _11491_ (.A(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__a22o_1 _11492_ (.A1(\r1.regblock[1][19] ),
    .A2(_06036_),
    .B1(_06037_),
    .B2(_06039_),
    .X(_02544_));
 sky130_fd_sc_hd__clkbuf_1 _11493_ (.A(_06033_),
    .X(_01518_));
 sky130_fd_sc_hd__buf_1 _11494_ (.A(_05669_),
    .X(_06040_));
 sky130_fd_sc_hd__a22o_1 _11495_ (.A1(\r1.regblock[1][18] ),
    .A2(_06036_),
    .B1(_06040_),
    .B2(_06039_),
    .X(_02543_));
 sky130_fd_sc_hd__buf_1 _11496_ (.A(_06032_),
    .X(_06041_));
 sky130_fd_sc_hd__buf_1 _11497_ (.A(_06041_),
    .X(_01517_));
 sky130_fd_sc_hd__buf_1 _11498_ (.A(_05673_),
    .X(_06042_));
 sky130_fd_sc_hd__a22o_1 _11499_ (.A1(\r1.regblock[1][17] ),
    .A2(_06036_),
    .B1(_06042_),
    .B2(_06039_),
    .X(_02542_));
 sky130_fd_sc_hd__clkbuf_1 _11500_ (.A(_06041_),
    .X(_01516_));
 sky130_fd_sc_hd__buf_1 _11501_ (.A(_06035_),
    .X(_06043_));
 sky130_fd_sc_hd__buf_1 _11502_ (.A(_05676_),
    .X(_06044_));
 sky130_fd_sc_hd__buf_1 _11503_ (.A(_06038_),
    .X(_06045_));
 sky130_fd_sc_hd__a22o_1 _11504_ (.A1(\r1.regblock[1][16] ),
    .A2(_06043_),
    .B1(_06044_),
    .B2(_06045_),
    .X(_02541_));
 sky130_fd_sc_hd__clkbuf_1 _11505_ (.A(_06041_),
    .X(_01515_));
 sky130_fd_sc_hd__buf_1 _11506_ (.A(_05679_),
    .X(_06046_));
 sky130_fd_sc_hd__a22o_1 _11507_ (.A1(\r1.regblock[1][15] ),
    .A2(_06043_),
    .B1(_06046_),
    .B2(_06045_),
    .X(_02540_));
 sky130_fd_sc_hd__buf_1 _11508_ (.A(_06032_),
    .X(_06047_));
 sky130_fd_sc_hd__clkbuf_1 _11509_ (.A(_06047_),
    .X(_01514_));
 sky130_fd_sc_hd__buf_1 _11510_ (.A(_05682_),
    .X(_06048_));
 sky130_fd_sc_hd__a22o_1 _11511_ (.A1(\r1.regblock[1][14] ),
    .A2(_06043_),
    .B1(_06048_),
    .B2(_06045_),
    .X(_02539_));
 sky130_fd_sc_hd__clkbuf_1 _11512_ (.A(_06047_),
    .X(_01513_));
 sky130_fd_sc_hd__buf_1 _11513_ (.A(_06035_),
    .X(_06049_));
 sky130_fd_sc_hd__buf_1 _11514_ (.A(_05685_),
    .X(_06050_));
 sky130_fd_sc_hd__buf_1 _11515_ (.A(_06038_),
    .X(_06051_));
 sky130_fd_sc_hd__a22o_1 _11516_ (.A1(\r1.regblock[1][13] ),
    .A2(_06049_),
    .B1(_06050_),
    .B2(_06051_),
    .X(_02538_));
 sky130_fd_sc_hd__clkbuf_1 _11517_ (.A(_06047_),
    .X(_01512_));
 sky130_fd_sc_hd__buf_1 _11518_ (.A(_05688_),
    .X(_06052_));
 sky130_fd_sc_hd__a22o_1 _11519_ (.A1(\r1.regblock[1][12] ),
    .A2(_06049_),
    .B1(_06052_),
    .B2(_06051_),
    .X(_02537_));
 sky130_fd_sc_hd__buf_1 _11520_ (.A(_06008_),
    .X(_06053_));
 sky130_fd_sc_hd__buf_1 _11521_ (.A(_06053_),
    .X(_06054_));
 sky130_fd_sc_hd__clkbuf_2 _11522_ (.A(_06054_),
    .X(_01511_));
 sky130_fd_sc_hd__buf_1 _11523_ (.A(_05691_),
    .X(_06055_));
 sky130_fd_sc_hd__a22o_1 _11524_ (.A1(\r1.regblock[1][11] ),
    .A2(_06049_),
    .B1(_06055_),
    .B2(_06051_),
    .X(_02536_));
 sky130_fd_sc_hd__clkbuf_1 _11525_ (.A(_06054_),
    .X(_01510_));
 sky130_fd_sc_hd__buf_1 _11526_ (.A(_06012_),
    .X(_06056_));
 sky130_fd_sc_hd__buf_1 _11527_ (.A(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__clkbuf_2 _11528_ (.A(_05695_),
    .X(_06058_));
 sky130_fd_sc_hd__buf_1 _11529_ (.A(_06016_),
    .X(_06059_));
 sky130_fd_sc_hd__buf_1 _11530_ (.A(_06059_),
    .X(_06060_));
 sky130_fd_sc_hd__a22o_1 _11531_ (.A1(\r1.regblock[1][10] ),
    .A2(_06057_),
    .B1(_06058_),
    .B2(_06060_),
    .X(_02535_));
 sky130_fd_sc_hd__clkbuf_1 _11532_ (.A(_06054_),
    .X(_01509_));
 sky130_fd_sc_hd__clkbuf_2 _11533_ (.A(_05699_),
    .X(_06061_));
 sky130_fd_sc_hd__a22o_1 _11534_ (.A1(\r1.regblock[1][9] ),
    .A2(_06057_),
    .B1(_06061_),
    .B2(_06060_),
    .X(_02534_));
 sky130_fd_sc_hd__buf_1 _11535_ (.A(_06053_),
    .X(_06062_));
 sky130_fd_sc_hd__clkbuf_1 _11536_ (.A(_06062_),
    .X(_01508_));
 sky130_fd_sc_hd__clkbuf_2 _11537_ (.A(_05703_),
    .X(_06063_));
 sky130_fd_sc_hd__a22o_1 _11538_ (.A1(\r1.regblock[1][8] ),
    .A2(_06057_),
    .B1(_06063_),
    .B2(_06060_),
    .X(_02533_));
 sky130_fd_sc_hd__clkbuf_1 _11539_ (.A(_06062_),
    .X(_01507_));
 sky130_fd_sc_hd__buf_1 _11540_ (.A(_06056_),
    .X(_06064_));
 sky130_fd_sc_hd__clkbuf_2 _11541_ (.A(_05706_),
    .X(_06065_));
 sky130_fd_sc_hd__buf_1 _11542_ (.A(_06059_),
    .X(_06066_));
 sky130_fd_sc_hd__a22o_1 _11543_ (.A1(\r1.regblock[1][7] ),
    .A2(_06064_),
    .B1(_06065_),
    .B2(_06066_),
    .X(_02532_));
 sky130_fd_sc_hd__clkbuf_1 _11544_ (.A(_06062_),
    .X(_01506_));
 sky130_fd_sc_hd__clkbuf_2 _11545_ (.A(_05709_),
    .X(_06067_));
 sky130_fd_sc_hd__a22o_1 _11546_ (.A1(\r1.regblock[1][6] ),
    .A2(_06064_),
    .B1(_06067_),
    .B2(_06066_),
    .X(_02531_));
 sky130_fd_sc_hd__buf_1 _11547_ (.A(_06053_),
    .X(_06068_));
 sky130_fd_sc_hd__clkbuf_1 _11548_ (.A(_06068_),
    .X(_01505_));
 sky130_fd_sc_hd__clkbuf_2 _11549_ (.A(_05712_),
    .X(_06069_));
 sky130_fd_sc_hd__a22o_1 _11550_ (.A1(\r1.regblock[1][5] ),
    .A2(_06064_),
    .B1(_06069_),
    .B2(_06066_),
    .X(_02530_));
 sky130_fd_sc_hd__clkbuf_1 _11551_ (.A(_06068_),
    .X(_01504_));
 sky130_fd_sc_hd__buf_1 _11552_ (.A(_06056_),
    .X(_06070_));
 sky130_fd_sc_hd__clkbuf_2 _11553_ (.A(_05715_),
    .X(_06071_));
 sky130_fd_sc_hd__buf_1 _11554_ (.A(_06059_),
    .X(_06072_));
 sky130_fd_sc_hd__a22o_1 _11555_ (.A1(\r1.regblock[1][4] ),
    .A2(_06070_),
    .B1(_06071_),
    .B2(_06072_),
    .X(_02529_));
 sky130_fd_sc_hd__clkbuf_1 _11556_ (.A(_06068_),
    .X(_01503_));
 sky130_fd_sc_hd__clkbuf_2 _11557_ (.A(_05718_),
    .X(_06073_));
 sky130_fd_sc_hd__a22o_1 _11558_ (.A1(\r1.regblock[1][3] ),
    .A2(_06070_),
    .B1(_06073_),
    .B2(_06072_),
    .X(_02528_));
 sky130_fd_sc_hd__buf_1 _11559_ (.A(_03907_),
    .X(_06074_));
 sky130_fd_sc_hd__buf_1 _11560_ (.A(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__buf_2 _11561_ (.A(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__buf_1 _11562_ (.A(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__buf_1 _11563_ (.A(_06077_),
    .X(_01502_));
 sky130_fd_sc_hd__clkbuf_2 _11564_ (.A(_05721_),
    .X(_06078_));
 sky130_fd_sc_hd__a22o_1 _11565_ (.A1(\r1.regblock[1][2] ),
    .A2(_06070_),
    .B1(_06078_),
    .B2(_06072_),
    .X(_02527_));
 sky130_fd_sc_hd__clkbuf_1 _11566_ (.A(_06077_),
    .X(_01501_));
 sky130_fd_sc_hd__buf_1 _11567_ (.A(_05723_),
    .X(_06079_));
 sky130_fd_sc_hd__a22o_1 _11568_ (.A1(\r1.regblock[1][1] ),
    .A2(_06001_),
    .B1(_06079_),
    .B2(_06005_),
    .X(_02526_));
 sky130_fd_sc_hd__clkbuf_1 _11569_ (.A(_06077_),
    .X(_01500_));
 sky130_fd_sc_hd__buf_1 _11570_ (.A(_05725_),
    .X(_06080_));
 sky130_fd_sc_hd__a22o_1 _11571_ (.A1(\r1.regblock[1][0] ),
    .A2(_06001_),
    .B1(_06080_),
    .B2(_06005_),
    .X(_02525_));
 sky130_fd_sc_hd__buf_1 _11572_ (.A(_06076_),
    .X(_06081_));
 sky130_fd_sc_hd__clkbuf_1 _11573_ (.A(_06081_),
    .X(_01499_));
 sky130_fd_sc_hd__or3_1 _11574_ (.A(_04340_),
    .B(_04214_),
    .C(_04392_),
    .X(_06082_));
 sky130_fd_sc_hd__clkbuf_1 _11575_ (.A(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__or2_2 _11576_ (.A(_04695_),
    .B(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__buf_1 _11577_ (.A(_06084_),
    .X(_06085_));
 sky130_fd_sc_hd__buf_1 _11578_ (.A(_06085_),
    .X(_06086_));
 sky130_fd_sc_hd__inv_2 _11579_ (.A(_06084_),
    .Y(_06087_));
 sky130_fd_sc_hd__buf_1 _11580_ (.A(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__buf_1 _11581_ (.A(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__a22o_1 _11582_ (.A1(\r1.regblock[20][31] ),
    .A2(_06086_),
    .B1(_06003_),
    .B2(_06089_),
    .X(_02524_));
 sky130_fd_sc_hd__clkbuf_1 _11583_ (.A(_06081_),
    .X(_01498_));
 sky130_fd_sc_hd__a22o_1 _11584_ (.A1(\r1.regblock[20][30] ),
    .A2(_06086_),
    .B1(_06007_),
    .B2(_06089_),
    .X(_02523_));
 sky130_fd_sc_hd__clkbuf_1 _11585_ (.A(_06081_),
    .X(_01497_));
 sky130_fd_sc_hd__a22o_1 _11586_ (.A1(\r1.regblock[20][29] ),
    .A2(_06086_),
    .B1(_06011_),
    .B2(_06089_),
    .X(_02522_));
 sky130_fd_sc_hd__buf_1 _11587_ (.A(_06076_),
    .X(_06090_));
 sky130_fd_sc_hd__clkbuf_1 _11588_ (.A(_06090_),
    .X(_01496_));
 sky130_fd_sc_hd__buf_2 _11589_ (.A(_06084_),
    .X(_06091_));
 sky130_fd_sc_hd__buf_2 _11590_ (.A(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__buf_1 _11591_ (.A(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__buf_2 _11592_ (.A(_06087_),
    .X(_06094_));
 sky130_fd_sc_hd__buf_2 _11593_ (.A(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__buf_1 _11594_ (.A(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__a22o_1 _11595_ (.A1(\r1.regblock[20][28] ),
    .A2(_06093_),
    .B1(_06015_),
    .B2(_06096_),
    .X(_02521_));
 sky130_fd_sc_hd__clkbuf_1 _11596_ (.A(_06090_),
    .X(_01495_));
 sky130_fd_sc_hd__a22o_1 _11597_ (.A1(\r1.regblock[20][27] ),
    .A2(_06093_),
    .B1(_06019_),
    .B2(_06096_),
    .X(_02520_));
 sky130_fd_sc_hd__clkbuf_1 _11598_ (.A(_06090_),
    .X(_01494_));
 sky130_fd_sc_hd__a22o_1 _11599_ (.A1(\r1.regblock[20][26] ),
    .A2(_06093_),
    .B1(_06021_),
    .B2(_06096_),
    .X(_02519_));
 sky130_fd_sc_hd__clkbuf_4 _11600_ (.A(_06075_),
    .X(_06097_));
 sky130_fd_sc_hd__buf_1 _11601_ (.A(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__clkbuf_1 _11602_ (.A(_06098_),
    .X(_01493_));
 sky130_fd_sc_hd__buf_1 _11603_ (.A(_06092_),
    .X(_06099_));
 sky130_fd_sc_hd__buf_1 _11604_ (.A(_06095_),
    .X(_06100_));
 sky130_fd_sc_hd__a22o_1 _11605_ (.A1(\r1.regblock[20][25] ),
    .A2(_06099_),
    .B1(_06023_),
    .B2(_06100_),
    .X(_02518_));
 sky130_fd_sc_hd__clkbuf_1 _11606_ (.A(_06098_),
    .X(_01492_));
 sky130_fd_sc_hd__a22o_1 _11607_ (.A1(\r1.regblock[20][24] ),
    .A2(_06099_),
    .B1(_06025_),
    .B2(_06100_),
    .X(_02517_));
 sky130_fd_sc_hd__clkbuf_1 _11608_ (.A(_06098_),
    .X(_01491_));
 sky130_fd_sc_hd__a22o_1 _11609_ (.A1(\r1.regblock[20][23] ),
    .A2(_06099_),
    .B1(_06027_),
    .B2(_06100_),
    .X(_02516_));
 sky130_fd_sc_hd__buf_1 _11610_ (.A(_06097_),
    .X(_06101_));
 sky130_fd_sc_hd__clkbuf_1 _11611_ (.A(_06101_),
    .X(_01490_));
 sky130_fd_sc_hd__buf_1 _11612_ (.A(_06092_),
    .X(_06102_));
 sky130_fd_sc_hd__buf_1 _11613_ (.A(_06095_),
    .X(_06103_));
 sky130_fd_sc_hd__a22o_1 _11614_ (.A1(\r1.regblock[20][22] ),
    .A2(_06102_),
    .B1(_06029_),
    .B2(_06103_),
    .X(_02515_));
 sky130_fd_sc_hd__clkbuf_1 _11615_ (.A(_06101_),
    .X(_01489_));
 sky130_fd_sc_hd__a22o_1 _11616_ (.A1(\r1.regblock[20][21] ),
    .A2(_06102_),
    .B1(_06031_),
    .B2(_06103_),
    .X(_02514_));
 sky130_fd_sc_hd__clkbuf_1 _11617_ (.A(_06101_),
    .X(_01488_));
 sky130_fd_sc_hd__a22o_1 _11618_ (.A1(\r1.regblock[20][20] ),
    .A2(_06102_),
    .B1(_06034_),
    .B2(_06103_),
    .X(_02513_));
 sky130_fd_sc_hd__buf_1 _11619_ (.A(_06097_),
    .X(_06104_));
 sky130_fd_sc_hd__clkbuf_1 _11620_ (.A(_06104_),
    .X(_01487_));
 sky130_fd_sc_hd__clkbuf_2 _11621_ (.A(_06091_),
    .X(_06105_));
 sky130_fd_sc_hd__buf_1 _11622_ (.A(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__clkbuf_2 _11623_ (.A(_06094_),
    .X(_06107_));
 sky130_fd_sc_hd__buf_1 _11624_ (.A(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__a22o_1 _11625_ (.A1(\r1.regblock[20][19] ),
    .A2(_06106_),
    .B1(_06037_),
    .B2(_06108_),
    .X(_02512_));
 sky130_fd_sc_hd__clkbuf_1 _11626_ (.A(_06104_),
    .X(_01486_));
 sky130_fd_sc_hd__a22o_1 _11627_ (.A1(\r1.regblock[20][18] ),
    .A2(_06106_),
    .B1(_06040_),
    .B2(_06108_),
    .X(_02511_));
 sky130_fd_sc_hd__clkbuf_1 _11628_ (.A(_06104_),
    .X(_01485_));
 sky130_fd_sc_hd__a22o_1 _11629_ (.A1(\r1.regblock[20][17] ),
    .A2(_06106_),
    .B1(_06042_),
    .B2(_06108_),
    .X(_02510_));
 sky130_fd_sc_hd__clkbuf_4 _11630_ (.A(_06075_),
    .X(_06109_));
 sky130_fd_sc_hd__buf_1 _11631_ (.A(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__clkbuf_1 _11632_ (.A(_06110_),
    .X(_01484_));
 sky130_fd_sc_hd__buf_1 _11633_ (.A(_06105_),
    .X(_06111_));
 sky130_fd_sc_hd__buf_1 _11634_ (.A(_06107_),
    .X(_06112_));
 sky130_fd_sc_hd__a22o_1 _11635_ (.A1(\r1.regblock[20][16] ),
    .A2(_06111_),
    .B1(_06044_),
    .B2(_06112_),
    .X(_02509_));
 sky130_fd_sc_hd__clkbuf_1 _11636_ (.A(_06110_),
    .X(_01483_));
 sky130_fd_sc_hd__a22o_1 _11637_ (.A1(\r1.regblock[20][15] ),
    .A2(_06111_),
    .B1(_06046_),
    .B2(_06112_),
    .X(_02508_));
 sky130_fd_sc_hd__clkbuf_1 _11638_ (.A(_06110_),
    .X(_01482_));
 sky130_fd_sc_hd__a22o_1 _11639_ (.A1(\r1.regblock[20][14] ),
    .A2(_06111_),
    .B1(_06048_),
    .B2(_06112_),
    .X(_02507_));
 sky130_fd_sc_hd__buf_1 _11640_ (.A(_06109_),
    .X(_06113_));
 sky130_fd_sc_hd__clkbuf_1 _11641_ (.A(_06113_),
    .X(_01481_));
 sky130_fd_sc_hd__buf_1 _11642_ (.A(_06105_),
    .X(_06114_));
 sky130_fd_sc_hd__buf_1 _11643_ (.A(_06107_),
    .X(_06115_));
 sky130_fd_sc_hd__a22o_1 _11644_ (.A1(\r1.regblock[20][13] ),
    .A2(_06114_),
    .B1(_06050_),
    .B2(_06115_),
    .X(_02506_));
 sky130_fd_sc_hd__clkbuf_1 _11645_ (.A(_06113_),
    .X(_01480_));
 sky130_fd_sc_hd__a22o_1 _11646_ (.A1(\r1.regblock[20][12] ),
    .A2(_06114_),
    .B1(_06052_),
    .B2(_06115_),
    .X(_02505_));
 sky130_fd_sc_hd__clkbuf_1 _11647_ (.A(_06113_),
    .X(_01479_));
 sky130_fd_sc_hd__a22o_1 _11648_ (.A1(\r1.regblock[20][11] ),
    .A2(_06114_),
    .B1(_06055_),
    .B2(_06115_),
    .X(_02504_));
 sky130_fd_sc_hd__buf_1 _11649_ (.A(_06109_),
    .X(_06116_));
 sky130_fd_sc_hd__clkbuf_1 _11650_ (.A(_06116_),
    .X(_01478_));
 sky130_fd_sc_hd__clkbuf_2 _11651_ (.A(_06091_),
    .X(_06117_));
 sky130_fd_sc_hd__buf_1 _11652_ (.A(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__clkbuf_2 _11653_ (.A(_06094_),
    .X(_06119_));
 sky130_fd_sc_hd__buf_1 _11654_ (.A(_06119_),
    .X(_06120_));
 sky130_fd_sc_hd__a22o_1 _11655_ (.A1(\r1.regblock[20][10] ),
    .A2(_06118_),
    .B1(_06058_),
    .B2(_06120_),
    .X(_02503_));
 sky130_fd_sc_hd__clkbuf_1 _11656_ (.A(_06116_),
    .X(_01477_));
 sky130_fd_sc_hd__a22o_1 _11657_ (.A1(\r1.regblock[20][9] ),
    .A2(_06118_),
    .B1(_06061_),
    .B2(_06120_),
    .X(_02502_));
 sky130_fd_sc_hd__clkbuf_1 _11658_ (.A(_06116_),
    .X(_01476_));
 sky130_fd_sc_hd__a22o_1 _11659_ (.A1(\r1.regblock[20][8] ),
    .A2(_06118_),
    .B1(_06063_),
    .B2(_06120_),
    .X(_02501_));
 sky130_fd_sc_hd__buf_1 _11660_ (.A(_06074_),
    .X(_06121_));
 sky130_fd_sc_hd__clkbuf_2 _11661_ (.A(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__buf_1 _11662_ (.A(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__clkbuf_1 _11663_ (.A(_06123_),
    .X(_01475_));
 sky130_fd_sc_hd__buf_1 _11664_ (.A(_06117_),
    .X(_06124_));
 sky130_fd_sc_hd__buf_1 _11665_ (.A(_06119_),
    .X(_06125_));
 sky130_fd_sc_hd__a22o_1 _11666_ (.A1(\r1.regblock[20][7] ),
    .A2(_06124_),
    .B1(_06065_),
    .B2(_06125_),
    .X(_02500_));
 sky130_fd_sc_hd__clkbuf_1 _11667_ (.A(_06123_),
    .X(_01474_));
 sky130_fd_sc_hd__a22o_1 _11668_ (.A1(\r1.regblock[20][6] ),
    .A2(_06124_),
    .B1(_06067_),
    .B2(_06125_),
    .X(_02499_));
 sky130_fd_sc_hd__clkbuf_1 _11669_ (.A(_06123_),
    .X(_01473_));
 sky130_fd_sc_hd__a22o_1 _11670_ (.A1(\r1.regblock[20][5] ),
    .A2(_06124_),
    .B1(_06069_),
    .B2(_06125_),
    .X(_02498_));
 sky130_fd_sc_hd__buf_1 _11671_ (.A(_06122_),
    .X(_06126_));
 sky130_fd_sc_hd__clkbuf_1 _11672_ (.A(_06126_),
    .X(_01472_));
 sky130_fd_sc_hd__buf_1 _11673_ (.A(_06117_),
    .X(_06127_));
 sky130_fd_sc_hd__buf_1 _11674_ (.A(_06119_),
    .X(_06128_));
 sky130_fd_sc_hd__a22o_1 _11675_ (.A1(\r1.regblock[20][4] ),
    .A2(_06127_),
    .B1(_06071_),
    .B2(_06128_),
    .X(_02497_));
 sky130_fd_sc_hd__clkbuf_1 _11676_ (.A(_06126_),
    .X(_01471_));
 sky130_fd_sc_hd__a22o_1 _11677_ (.A1(\r1.regblock[20][3] ),
    .A2(_06127_),
    .B1(_06073_),
    .B2(_06128_),
    .X(_02496_));
 sky130_fd_sc_hd__clkbuf_1 _11678_ (.A(_06126_),
    .X(_01470_));
 sky130_fd_sc_hd__a22o_1 _11679_ (.A1(\r1.regblock[20][2] ),
    .A2(_06127_),
    .B1(_06078_),
    .B2(_06128_),
    .X(_02495_));
 sky130_fd_sc_hd__buf_1 _11680_ (.A(_06122_),
    .X(_06129_));
 sky130_fd_sc_hd__clkbuf_1 _11681_ (.A(_06129_),
    .X(_01469_));
 sky130_fd_sc_hd__a22o_1 _11682_ (.A1(\r1.regblock[20][1] ),
    .A2(_06085_),
    .B1(_06079_),
    .B2(_06088_),
    .X(_02494_));
 sky130_fd_sc_hd__clkbuf_1 _11683_ (.A(_06129_),
    .X(_01468_));
 sky130_fd_sc_hd__a22o_1 _11684_ (.A1(\r1.regblock[20][0] ),
    .A2(_06085_),
    .B1(_06080_),
    .B2(_06088_),
    .X(_02493_));
 sky130_fd_sc_hd__clkbuf_1 _11685_ (.A(_06129_),
    .X(_01467_));
 sky130_fd_sc_hd__or2_2 _11686_ (.A(_04396_),
    .B(_06083_),
    .X(_06130_));
 sky130_fd_sc_hd__buf_1 _11687_ (.A(_06130_),
    .X(_06131_));
 sky130_fd_sc_hd__buf_1 _11688_ (.A(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__inv_2 _11689_ (.A(_06130_),
    .Y(_06133_));
 sky130_fd_sc_hd__buf_1 _11690_ (.A(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__buf_1 _11691_ (.A(_06134_),
    .X(_06135_));
 sky130_fd_sc_hd__a22o_1 _11692_ (.A1(\r1.regblock[21][31] ),
    .A2(_06132_),
    .B1(_06003_),
    .B2(_06135_),
    .X(_02492_));
 sky130_fd_sc_hd__buf_2 _11693_ (.A(_06121_),
    .X(_06136_));
 sky130_fd_sc_hd__buf_1 _11694_ (.A(_06136_),
    .X(_06137_));
 sky130_fd_sc_hd__clkbuf_1 _11695_ (.A(_06137_),
    .X(_01466_));
 sky130_fd_sc_hd__a22o_1 _11696_ (.A1(\r1.regblock[21][30] ),
    .A2(_06132_),
    .B1(_06007_),
    .B2(_06135_),
    .X(_02491_));
 sky130_fd_sc_hd__clkbuf_1 _11697_ (.A(_06137_),
    .X(_01465_));
 sky130_fd_sc_hd__a22o_1 _11698_ (.A1(\r1.regblock[21][29] ),
    .A2(_06132_),
    .B1(_06011_),
    .B2(_06135_),
    .X(_02490_));
 sky130_fd_sc_hd__clkbuf_1 _11699_ (.A(_06137_),
    .X(_01464_));
 sky130_fd_sc_hd__clkbuf_2 _11700_ (.A(_06130_),
    .X(_06138_));
 sky130_fd_sc_hd__buf_2 _11701_ (.A(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__buf_1 _11702_ (.A(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__buf_2 _11703_ (.A(_06133_),
    .X(_06141_));
 sky130_fd_sc_hd__buf_2 _11704_ (.A(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__buf_1 _11705_ (.A(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__a22o_1 _11706_ (.A1(\r1.regblock[21][28] ),
    .A2(_06140_),
    .B1(_06015_),
    .B2(_06143_),
    .X(_02489_));
 sky130_fd_sc_hd__buf_1 _11707_ (.A(_06136_),
    .X(_06144_));
 sky130_fd_sc_hd__clkbuf_1 _11708_ (.A(_06144_),
    .X(_01463_));
 sky130_fd_sc_hd__a22o_1 _11709_ (.A1(\r1.regblock[21][27] ),
    .A2(_06140_),
    .B1(_06019_),
    .B2(_06143_),
    .X(_02488_));
 sky130_fd_sc_hd__clkbuf_1 _11710_ (.A(_06144_),
    .X(_01462_));
 sky130_fd_sc_hd__a22o_1 _11711_ (.A1(\r1.regblock[21][26] ),
    .A2(_06140_),
    .B1(_06021_),
    .B2(_06143_),
    .X(_02487_));
 sky130_fd_sc_hd__clkbuf_1 _11712_ (.A(_06144_),
    .X(_01461_));
 sky130_fd_sc_hd__buf_1 _11713_ (.A(_06139_),
    .X(_06145_));
 sky130_fd_sc_hd__buf_1 _11714_ (.A(_06142_),
    .X(_06146_));
 sky130_fd_sc_hd__a22o_1 _11715_ (.A1(\r1.regblock[21][25] ),
    .A2(_06145_),
    .B1(_06023_),
    .B2(_06146_),
    .X(_02486_));
 sky130_fd_sc_hd__clkbuf_2 _11716_ (.A(_06136_),
    .X(_06147_));
 sky130_fd_sc_hd__clkbuf_1 _11717_ (.A(_06147_),
    .X(_01460_));
 sky130_fd_sc_hd__a22o_1 _11718_ (.A1(\r1.regblock[21][24] ),
    .A2(_06145_),
    .B1(_06025_),
    .B2(_06146_),
    .X(_02485_));
 sky130_fd_sc_hd__clkbuf_1 _11719_ (.A(_06147_),
    .X(_01459_));
 sky130_fd_sc_hd__a22o_1 _11720_ (.A1(\r1.regblock[21][23] ),
    .A2(_06145_),
    .B1(_06027_),
    .B2(_06146_),
    .X(_02484_));
 sky130_fd_sc_hd__clkbuf_1 _11721_ (.A(_06147_),
    .X(_01458_));
 sky130_fd_sc_hd__buf_1 _11722_ (.A(_06139_),
    .X(_06148_));
 sky130_fd_sc_hd__buf_1 _11723_ (.A(_06142_),
    .X(_06149_));
 sky130_fd_sc_hd__a22o_1 _11724_ (.A1(\r1.regblock[21][22] ),
    .A2(_06148_),
    .B1(_06029_),
    .B2(_06149_),
    .X(_02483_));
 sky130_fd_sc_hd__clkbuf_2 _11725_ (.A(_06121_),
    .X(_06150_));
 sky130_fd_sc_hd__clkbuf_2 _11726_ (.A(_06150_),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_1 _11727_ (.A(_06151_),
    .X(_01457_));
 sky130_fd_sc_hd__a22o_1 _11728_ (.A1(\r1.regblock[21][21] ),
    .A2(_06148_),
    .B1(_06031_),
    .B2(_06149_),
    .X(_02482_));
 sky130_fd_sc_hd__clkbuf_1 _11729_ (.A(_06151_),
    .X(_01456_));
 sky130_fd_sc_hd__a22o_1 _11730_ (.A1(\r1.regblock[21][20] ),
    .A2(_06148_),
    .B1(_06034_),
    .B2(_06149_),
    .X(_02481_));
 sky130_fd_sc_hd__clkbuf_1 _11731_ (.A(_06151_),
    .X(_01455_));
 sky130_fd_sc_hd__clkbuf_2 _11732_ (.A(_06138_),
    .X(_06152_));
 sky130_fd_sc_hd__buf_1 _11733_ (.A(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__clkbuf_2 _11734_ (.A(_06141_),
    .X(_06154_));
 sky130_fd_sc_hd__buf_1 _11735_ (.A(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__a22o_1 _11736_ (.A1(\r1.regblock[21][19] ),
    .A2(_06153_),
    .B1(_06037_),
    .B2(_06155_),
    .X(_02480_));
 sky130_fd_sc_hd__buf_1 _11737_ (.A(_06150_),
    .X(_06156_));
 sky130_fd_sc_hd__clkbuf_1 _11738_ (.A(_06156_),
    .X(_01454_));
 sky130_fd_sc_hd__a22o_1 _11739_ (.A1(\r1.regblock[21][18] ),
    .A2(_06153_),
    .B1(_06040_),
    .B2(_06155_),
    .X(_02479_));
 sky130_fd_sc_hd__clkbuf_1 _11740_ (.A(_06156_),
    .X(_01453_));
 sky130_fd_sc_hd__a22o_1 _11741_ (.A1(\r1.regblock[21][17] ),
    .A2(_06153_),
    .B1(_06042_),
    .B2(_06155_),
    .X(_02478_));
 sky130_fd_sc_hd__clkbuf_1 _11742_ (.A(_06156_),
    .X(_01452_));
 sky130_fd_sc_hd__buf_1 _11743_ (.A(_06152_),
    .X(_06157_));
 sky130_fd_sc_hd__buf_1 _11744_ (.A(_06154_),
    .X(_06158_));
 sky130_fd_sc_hd__a22o_1 _11745_ (.A1(\r1.regblock[21][16] ),
    .A2(_06157_),
    .B1(_06044_),
    .B2(_06158_),
    .X(_02477_));
 sky130_fd_sc_hd__buf_1 _11746_ (.A(_06150_),
    .X(_06159_));
 sky130_fd_sc_hd__clkbuf_1 _11747_ (.A(_06159_),
    .X(_01451_));
 sky130_fd_sc_hd__a22o_1 _11748_ (.A1(\r1.regblock[21][15] ),
    .A2(_06157_),
    .B1(_06046_),
    .B2(_06158_),
    .X(_02476_));
 sky130_fd_sc_hd__clkbuf_1 _11749_ (.A(_06159_),
    .X(_01450_));
 sky130_fd_sc_hd__a22o_1 _11750_ (.A1(\r1.regblock[21][14] ),
    .A2(_06157_),
    .B1(_06048_),
    .B2(_06158_),
    .X(_02475_));
 sky130_fd_sc_hd__buf_1 _11751_ (.A(_06159_),
    .X(_01449_));
 sky130_fd_sc_hd__clkbuf_2 _11752_ (.A(_06152_),
    .X(_06160_));
 sky130_fd_sc_hd__buf_1 _11753_ (.A(_06154_),
    .X(_06161_));
 sky130_fd_sc_hd__a22o_1 _11754_ (.A1(\r1.regblock[21][13] ),
    .A2(_06160_),
    .B1(_06050_),
    .B2(_06161_),
    .X(_02474_));
 sky130_fd_sc_hd__clkbuf_2 _11755_ (.A(_06074_),
    .X(_06162_));
 sky130_fd_sc_hd__clkbuf_2 _11756_ (.A(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__clkbuf_2 _11757_ (.A(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__clkbuf_1 _11758_ (.A(_06164_),
    .X(_01448_));
 sky130_fd_sc_hd__a22o_1 _11759_ (.A1(\r1.regblock[21][12] ),
    .A2(_06160_),
    .B1(_06052_),
    .B2(_06161_),
    .X(_02473_));
 sky130_fd_sc_hd__clkbuf_1 _11760_ (.A(_06164_),
    .X(_01447_));
 sky130_fd_sc_hd__a22o_1 _11761_ (.A1(\r1.regblock[21][11] ),
    .A2(_06160_),
    .B1(_06055_),
    .B2(_06161_),
    .X(_02472_));
 sky130_fd_sc_hd__clkbuf_1 _11762_ (.A(_06164_),
    .X(_01446_));
 sky130_fd_sc_hd__buf_1 _11763_ (.A(_06138_),
    .X(_06165_));
 sky130_fd_sc_hd__buf_1 _11764_ (.A(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__buf_1 _11765_ (.A(_06141_),
    .X(_06167_));
 sky130_fd_sc_hd__buf_1 _11766_ (.A(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__a22o_1 _11767_ (.A1(\r1.regblock[21][10] ),
    .A2(_06166_),
    .B1(_06058_),
    .B2(_06168_),
    .X(_02471_));
 sky130_fd_sc_hd__buf_1 _11768_ (.A(_06163_),
    .X(_06169_));
 sky130_fd_sc_hd__clkbuf_1 _11769_ (.A(_06169_),
    .X(_01445_));
 sky130_fd_sc_hd__a22o_1 _11770_ (.A1(\r1.regblock[21][9] ),
    .A2(_06166_),
    .B1(_06061_),
    .B2(_06168_),
    .X(_02470_));
 sky130_fd_sc_hd__clkbuf_1 _11771_ (.A(_06169_),
    .X(_01444_));
 sky130_fd_sc_hd__a22o_1 _11772_ (.A1(\r1.regblock[21][8] ),
    .A2(_06166_),
    .B1(_06063_),
    .B2(_06168_),
    .X(_02469_));
 sky130_fd_sc_hd__clkbuf_1 _11773_ (.A(_06169_),
    .X(_01443_));
 sky130_fd_sc_hd__buf_1 _11774_ (.A(_06165_),
    .X(_06170_));
 sky130_fd_sc_hd__buf_1 _11775_ (.A(_06167_),
    .X(_06171_));
 sky130_fd_sc_hd__a22o_1 _11776_ (.A1(\r1.regblock[21][7] ),
    .A2(_06170_),
    .B1(_06065_),
    .B2(_06171_),
    .X(_02468_));
 sky130_fd_sc_hd__buf_1 _11777_ (.A(_06163_),
    .X(_06172_));
 sky130_fd_sc_hd__clkbuf_1 _11778_ (.A(_06172_),
    .X(_01442_));
 sky130_fd_sc_hd__a22o_1 _11779_ (.A1(\r1.regblock[21][6] ),
    .A2(_06170_),
    .B1(_06067_),
    .B2(_06171_),
    .X(_02467_));
 sky130_fd_sc_hd__clkbuf_1 _11780_ (.A(_06172_),
    .X(_01441_));
 sky130_fd_sc_hd__a22o_1 _11781_ (.A1(\r1.regblock[21][5] ),
    .A2(_06170_),
    .B1(_06069_),
    .B2(_06171_),
    .X(_02466_));
 sky130_fd_sc_hd__clkbuf_1 _11782_ (.A(_06172_),
    .X(_01440_));
 sky130_fd_sc_hd__buf_1 _11783_ (.A(_06165_),
    .X(_06173_));
 sky130_fd_sc_hd__buf_1 _11784_ (.A(_06167_),
    .X(_06174_));
 sky130_fd_sc_hd__a22o_1 _11785_ (.A1(\r1.regblock[21][4] ),
    .A2(_06173_),
    .B1(_06071_),
    .B2(_06174_),
    .X(_02465_));
 sky130_fd_sc_hd__buf_1 _11786_ (.A(_06162_),
    .X(_06175_));
 sky130_fd_sc_hd__clkbuf_2 _11787_ (.A(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__clkbuf_1 _11788_ (.A(_06176_),
    .X(_01439_));
 sky130_fd_sc_hd__a22o_1 _11789_ (.A1(\r1.regblock[21][3] ),
    .A2(_06173_),
    .B1(_06073_),
    .B2(_06174_),
    .X(_02464_));
 sky130_fd_sc_hd__clkbuf_1 _11790_ (.A(_06176_),
    .X(_01438_));
 sky130_fd_sc_hd__a22o_1 _11791_ (.A1(\r1.regblock[21][2] ),
    .A2(_06173_),
    .B1(_06078_),
    .B2(_06174_),
    .X(_02463_));
 sky130_fd_sc_hd__clkbuf_1 _11792_ (.A(_06176_),
    .X(_01437_));
 sky130_fd_sc_hd__a22o_1 _11793_ (.A1(\r1.regblock[21][1] ),
    .A2(_06131_),
    .B1(_06079_),
    .B2(_06134_),
    .X(_02462_));
 sky130_fd_sc_hd__buf_1 _11794_ (.A(_06175_),
    .X(_06177_));
 sky130_fd_sc_hd__clkbuf_1 _11795_ (.A(_06177_),
    .X(_01436_));
 sky130_fd_sc_hd__a22o_1 _11796_ (.A1(\r1.regblock[21][0] ),
    .A2(_06131_),
    .B1(_06080_),
    .B2(_06134_),
    .X(_02461_));
 sky130_fd_sc_hd__clkbuf_1 _11797_ (.A(_06177_),
    .X(_01435_));
 sky130_fd_sc_hd__or2_2 _11798_ (.A(_04449_),
    .B(_06083_),
    .X(_06178_));
 sky130_fd_sc_hd__buf_1 _11799_ (.A(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__buf_1 _11800_ (.A(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__inv_2 _11801_ (.A(_06178_),
    .Y(_06181_));
 sky130_fd_sc_hd__buf_1 _11802_ (.A(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__buf_1 _11803_ (.A(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__a22o_1 _11804_ (.A1(\r1.regblock[22][31] ),
    .A2(_06180_),
    .B1(_04228_),
    .B2(_06183_),
    .X(_02460_));
 sky130_fd_sc_hd__clkbuf_1 _11805_ (.A(_06177_),
    .X(_01434_));
 sky130_fd_sc_hd__a22o_1 _11806_ (.A1(\r1.regblock[22][30] ),
    .A2(_06180_),
    .B1(_04233_),
    .B2(_06183_),
    .X(_02459_));
 sky130_fd_sc_hd__clkbuf_2 _11807_ (.A(_06175_),
    .X(_06184_));
 sky130_fd_sc_hd__clkbuf_1 _11808_ (.A(_06184_),
    .X(_01433_));
 sky130_fd_sc_hd__a22o_1 _11809_ (.A1(\r1.regblock[22][29] ),
    .A2(_06180_),
    .B1(_04239_),
    .B2(_06183_),
    .X(_02458_));
 sky130_fd_sc_hd__clkbuf_1 _11810_ (.A(_06184_),
    .X(_01432_));
 sky130_fd_sc_hd__clkbuf_2 _11811_ (.A(_06178_),
    .X(_06185_));
 sky130_fd_sc_hd__buf_2 _11812_ (.A(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__buf_1 _11813_ (.A(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__clkbuf_2 _11814_ (.A(_06181_),
    .X(_06188_));
 sky130_fd_sc_hd__buf_2 _11815_ (.A(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__buf_1 _11816_ (.A(_06189_),
    .X(_06190_));
 sky130_fd_sc_hd__a22o_1 _11817_ (.A1(\r1.regblock[22][28] ),
    .A2(_06187_),
    .B1(_04244_),
    .B2(_06190_),
    .X(_02457_));
 sky130_fd_sc_hd__clkbuf_1 _11818_ (.A(_06184_),
    .X(_01431_));
 sky130_fd_sc_hd__a22o_1 _11819_ (.A1(\r1.regblock[22][27] ),
    .A2(_06187_),
    .B1(_04249_),
    .B2(_06190_),
    .X(_02456_));
 sky130_fd_sc_hd__clkbuf_2 _11820_ (.A(_06162_),
    .X(_06191_));
 sky130_fd_sc_hd__buf_1 _11821_ (.A(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__clkbuf_1 _11822_ (.A(_06192_),
    .X(_01430_));
 sky130_fd_sc_hd__a22o_1 _11823_ (.A1(\r1.regblock[22][26] ),
    .A2(_06187_),
    .B1(_04252_),
    .B2(_06190_),
    .X(_02455_));
 sky130_fd_sc_hd__clkbuf_1 _11824_ (.A(_06192_),
    .X(_01429_));
 sky130_fd_sc_hd__buf_1 _11825_ (.A(_06186_),
    .X(_06193_));
 sky130_fd_sc_hd__buf_1 _11826_ (.A(_06189_),
    .X(_06194_));
 sky130_fd_sc_hd__a22o_1 _11827_ (.A1(\r1.regblock[22][25] ),
    .A2(_06193_),
    .B1(_04255_),
    .B2(_06194_),
    .X(_02454_));
 sky130_fd_sc_hd__clkbuf_1 _11828_ (.A(_06192_),
    .X(_01428_));
 sky130_fd_sc_hd__a22o_1 _11829_ (.A1(\r1.regblock[22][24] ),
    .A2(_06193_),
    .B1(_04258_),
    .B2(_06194_),
    .X(_02453_));
 sky130_fd_sc_hd__clkbuf_2 _11830_ (.A(_06191_),
    .X(_06195_));
 sky130_fd_sc_hd__clkbuf_1 _11831_ (.A(_06195_),
    .X(_01427_));
 sky130_fd_sc_hd__a22o_1 _11832_ (.A1(\r1.regblock[22][23] ),
    .A2(_06193_),
    .B1(_04261_),
    .B2(_06194_),
    .X(_02452_));
 sky130_fd_sc_hd__clkbuf_1 _11833_ (.A(_06195_),
    .X(_01426_));
 sky130_fd_sc_hd__buf_1 _11834_ (.A(_06186_),
    .X(_06196_));
 sky130_fd_sc_hd__buf_1 _11835_ (.A(_06189_),
    .X(_06197_));
 sky130_fd_sc_hd__a22o_1 _11836_ (.A1(\r1.regblock[22][22] ),
    .A2(_06196_),
    .B1(_04264_),
    .B2(_06197_),
    .X(_02451_));
 sky130_fd_sc_hd__clkbuf_1 _11837_ (.A(_06195_),
    .X(_01425_));
 sky130_fd_sc_hd__a22o_1 _11838_ (.A1(\r1.regblock[22][21] ),
    .A2(_06196_),
    .B1(_04267_),
    .B2(_06197_),
    .X(_02450_));
 sky130_fd_sc_hd__clkbuf_2 _11839_ (.A(_06191_),
    .X(_06198_));
 sky130_fd_sc_hd__clkbuf_1 _11840_ (.A(_06198_),
    .X(_01424_));
 sky130_fd_sc_hd__a22o_1 _11841_ (.A1(\r1.regblock[22][20] ),
    .A2(_06196_),
    .B1(_04271_),
    .B2(_06197_),
    .X(_02449_));
 sky130_fd_sc_hd__clkbuf_1 _11842_ (.A(_06198_),
    .X(_01423_));
 sky130_fd_sc_hd__clkbuf_2 _11843_ (.A(_06185_),
    .X(_06199_));
 sky130_fd_sc_hd__buf_1 _11844_ (.A(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__clkbuf_2 _11845_ (.A(_06188_),
    .X(_06201_));
 sky130_fd_sc_hd__buf_1 _11846_ (.A(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__a22o_1 _11847_ (.A1(\r1.regblock[22][19] ),
    .A2(_06200_),
    .B1(_04275_),
    .B2(_06202_),
    .X(_02448_));
 sky130_fd_sc_hd__clkbuf_1 _11848_ (.A(_06198_),
    .X(_01422_));
 sky130_fd_sc_hd__a22o_1 _11849_ (.A1(\r1.regblock[22][18] ),
    .A2(_06200_),
    .B1(_04279_),
    .B2(_06202_),
    .X(_02447_));
 sky130_fd_sc_hd__buf_1 _11850_ (.A(_03908_),
    .X(_06203_));
 sky130_fd_sc_hd__clkbuf_4 _11851_ (.A(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__buf_1 _11852_ (.A(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__buf_1 _11853_ (.A(_06205_),
    .X(_01421_));
 sky130_fd_sc_hd__a22o_1 _11854_ (.A1(\r1.regblock[22][17] ),
    .A2(_06200_),
    .B1(_04282_),
    .B2(_06202_),
    .X(_02446_));
 sky130_fd_sc_hd__clkbuf_1 _11855_ (.A(_06205_),
    .X(_01420_));
 sky130_fd_sc_hd__buf_1 _11856_ (.A(_06199_),
    .X(_06206_));
 sky130_fd_sc_hd__buf_1 _11857_ (.A(_06201_),
    .X(_06207_));
 sky130_fd_sc_hd__a22o_1 _11858_ (.A1(\r1.regblock[22][16] ),
    .A2(_06206_),
    .B1(_04285_),
    .B2(_06207_),
    .X(_02445_));
 sky130_fd_sc_hd__clkbuf_1 _11859_ (.A(_06205_),
    .X(_01419_));
 sky130_fd_sc_hd__a22o_1 _11860_ (.A1(\r1.regblock[22][15] ),
    .A2(_06206_),
    .B1(_04288_),
    .B2(_06207_),
    .X(_02444_));
 sky130_fd_sc_hd__buf_1 _11861_ (.A(_06204_),
    .X(_06208_));
 sky130_fd_sc_hd__clkbuf_1 _11862_ (.A(_06208_),
    .X(_01418_));
 sky130_fd_sc_hd__a22o_1 _11863_ (.A1(\r1.regblock[22][14] ),
    .A2(_06206_),
    .B1(_04291_),
    .B2(_06207_),
    .X(_02443_));
 sky130_fd_sc_hd__clkbuf_1 _11864_ (.A(_06208_),
    .X(_01417_));
 sky130_fd_sc_hd__buf_1 _11865_ (.A(_06199_),
    .X(_06209_));
 sky130_fd_sc_hd__buf_1 _11866_ (.A(_06201_),
    .X(_06210_));
 sky130_fd_sc_hd__a22o_1 _11867_ (.A1(\r1.regblock[22][13] ),
    .A2(_06209_),
    .B1(_04294_),
    .B2(_06210_),
    .X(_02442_));
 sky130_fd_sc_hd__clkbuf_1 _11868_ (.A(_06208_),
    .X(_01416_));
 sky130_fd_sc_hd__a22o_1 _11869_ (.A1(\r1.regblock[22][12] ),
    .A2(_06209_),
    .B1(_04297_),
    .B2(_06210_),
    .X(_02441_));
 sky130_fd_sc_hd__buf_2 _11870_ (.A(_06204_),
    .X(_06211_));
 sky130_fd_sc_hd__clkbuf_1 _11871_ (.A(_06211_),
    .X(_01415_));
 sky130_fd_sc_hd__a22o_1 _11872_ (.A1(\r1.regblock[22][11] ),
    .A2(_06209_),
    .B1(_04301_),
    .B2(_06210_),
    .X(_02440_));
 sky130_fd_sc_hd__clkbuf_1 _11873_ (.A(_06211_),
    .X(_01414_));
 sky130_fd_sc_hd__clkbuf_2 _11874_ (.A(_06185_),
    .X(_06212_));
 sky130_fd_sc_hd__buf_1 _11875_ (.A(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__clkbuf_2 _11876_ (.A(_06188_),
    .X(_06214_));
 sky130_fd_sc_hd__buf_1 _11877_ (.A(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__a22o_1 _11878_ (.A1(\r1.regblock[22][10] ),
    .A2(_06213_),
    .B1(_04305_),
    .B2(_06215_),
    .X(_02439_));
 sky130_fd_sc_hd__clkbuf_1 _11879_ (.A(_06211_),
    .X(_01413_));
 sky130_fd_sc_hd__a22o_1 _11880_ (.A1(\r1.regblock[22][9] ),
    .A2(_06213_),
    .B1(_04309_),
    .B2(_06215_),
    .X(_02438_));
 sky130_fd_sc_hd__buf_1 _11881_ (.A(_06203_),
    .X(_06216_));
 sky130_fd_sc_hd__buf_1 _11882_ (.A(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__clkbuf_1 _11883_ (.A(_06217_),
    .X(_01412_));
 sky130_fd_sc_hd__a22o_1 _11884_ (.A1(\r1.regblock[22][8] ),
    .A2(_06213_),
    .B1(_04312_),
    .B2(_06215_),
    .X(_02437_));
 sky130_fd_sc_hd__clkbuf_1 _11885_ (.A(_06217_),
    .X(_01411_));
 sky130_fd_sc_hd__buf_1 _11886_ (.A(_06212_),
    .X(_06218_));
 sky130_fd_sc_hd__buf_1 _11887_ (.A(_06214_),
    .X(_06219_));
 sky130_fd_sc_hd__a22o_1 _11888_ (.A1(\r1.regblock[22][7] ),
    .A2(_06218_),
    .B1(_04315_),
    .B2(_06219_),
    .X(_02436_));
 sky130_fd_sc_hd__clkbuf_1 _11889_ (.A(_06217_),
    .X(_01410_));
 sky130_fd_sc_hd__a22o_1 _11890_ (.A1(\r1.regblock[22][6] ),
    .A2(_06218_),
    .B1(_04318_),
    .B2(_06219_),
    .X(_02435_));
 sky130_fd_sc_hd__buf_1 _11891_ (.A(_06216_),
    .X(_06220_));
 sky130_fd_sc_hd__clkbuf_1 _11892_ (.A(_06220_),
    .X(_01409_));
 sky130_fd_sc_hd__a22o_1 _11893_ (.A1(\r1.regblock[22][5] ),
    .A2(_06218_),
    .B1(_04321_),
    .B2(_06219_),
    .X(_02434_));
 sky130_fd_sc_hd__clkbuf_1 _11894_ (.A(_06220_),
    .X(_01408_));
 sky130_fd_sc_hd__buf_1 _11895_ (.A(_06212_),
    .X(_06221_));
 sky130_fd_sc_hd__buf_1 _11896_ (.A(_06214_),
    .X(_06222_));
 sky130_fd_sc_hd__a22o_1 _11897_ (.A1(\r1.regblock[22][4] ),
    .A2(_06221_),
    .B1(_04324_),
    .B2(_06222_),
    .X(_02433_));
 sky130_fd_sc_hd__clkbuf_1 _11898_ (.A(_06220_),
    .X(_01407_));
 sky130_fd_sc_hd__a22o_1 _11899_ (.A1(\r1.regblock[22][3] ),
    .A2(_06221_),
    .B1(_04327_),
    .B2(_06222_),
    .X(_02432_));
 sky130_fd_sc_hd__clkbuf_2 _11900_ (.A(_06216_),
    .X(_06223_));
 sky130_fd_sc_hd__clkbuf_1 _11901_ (.A(_06223_),
    .X(_01406_));
 sky130_fd_sc_hd__a22o_1 _11902_ (.A1(\r1.regblock[22][2] ),
    .A2(_06221_),
    .B1(_04332_),
    .B2(_06222_),
    .X(_02431_));
 sky130_fd_sc_hd__clkbuf_1 _11903_ (.A(_06223_),
    .X(_01405_));
 sky130_fd_sc_hd__a22o_1 _11904_ (.A1(\r1.regblock[22][1] ),
    .A2(_06179_),
    .B1(_04334_),
    .B2(_06182_),
    .X(_02430_));
 sky130_fd_sc_hd__clkbuf_1 _11905_ (.A(_06223_),
    .X(_01404_));
 sky130_fd_sc_hd__a22o_1 _11906_ (.A1(\r1.regblock[22][0] ),
    .A2(_06179_),
    .B1(_04336_),
    .B2(_06182_),
    .X(_02429_));
 sky130_fd_sc_hd__buf_2 _11907_ (.A(_06203_),
    .X(_06224_));
 sky130_fd_sc_hd__buf_1 _11908_ (.A(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__clkbuf_1 _11909_ (.A(_06225_),
    .X(_01403_));
 sky130_fd_sc_hd__or2_2 _11910_ (.A(_04224_),
    .B(_06082_),
    .X(_06226_));
 sky130_fd_sc_hd__buf_1 _11911_ (.A(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__buf_1 _11912_ (.A(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__inv_2 _11913_ (.A(_06226_),
    .Y(_06229_));
 sky130_fd_sc_hd__buf_1 _11914_ (.A(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__buf_1 _11915_ (.A(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__a22o_1 _11916_ (.A1(\r1.regblock[23][31] ),
    .A2(_06228_),
    .B1(_04228_),
    .B2(_06231_),
    .X(_02428_));
 sky130_fd_sc_hd__clkbuf_1 _11917_ (.A(_06225_),
    .X(_01402_));
 sky130_fd_sc_hd__a22o_1 _11918_ (.A1(\r1.regblock[23][30] ),
    .A2(_06228_),
    .B1(_04233_),
    .B2(_06231_),
    .X(_02427_));
 sky130_fd_sc_hd__clkbuf_1 _11919_ (.A(_06225_),
    .X(_01401_));
 sky130_fd_sc_hd__a22o_1 _11920_ (.A1(\r1.regblock[23][29] ),
    .A2(_06228_),
    .B1(_04239_),
    .B2(_06231_),
    .X(_02426_));
 sky130_fd_sc_hd__buf_1 _11921_ (.A(_06224_),
    .X(_06232_));
 sky130_fd_sc_hd__clkbuf_1 _11922_ (.A(_06232_),
    .X(_01400_));
 sky130_fd_sc_hd__clkbuf_2 _11923_ (.A(_06226_),
    .X(_06233_));
 sky130_fd_sc_hd__buf_2 _11924_ (.A(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__buf_1 _11925_ (.A(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__buf_2 _11926_ (.A(_06229_),
    .X(_06236_));
 sky130_fd_sc_hd__buf_2 _11927_ (.A(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__buf_1 _11928_ (.A(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__a22o_1 _11929_ (.A1(\r1.regblock[23][28] ),
    .A2(_06235_),
    .B1(_04244_),
    .B2(_06238_),
    .X(_02425_));
 sky130_fd_sc_hd__clkbuf_1 _11930_ (.A(_06232_),
    .X(_01399_));
 sky130_fd_sc_hd__a22o_1 _11931_ (.A1(\r1.regblock[23][27] ),
    .A2(_06235_),
    .B1(_04249_),
    .B2(_06238_),
    .X(_02424_));
 sky130_fd_sc_hd__clkbuf_1 _11932_ (.A(_06232_),
    .X(_01398_));
 sky130_fd_sc_hd__a22o_1 _11933_ (.A1(\r1.regblock[23][26] ),
    .A2(_06235_),
    .B1(_04252_),
    .B2(_06238_),
    .X(_02423_));
 sky130_fd_sc_hd__buf_1 _11934_ (.A(_06224_),
    .X(_06239_));
 sky130_fd_sc_hd__clkbuf_1 _11935_ (.A(_06239_),
    .X(_01397_));
 sky130_fd_sc_hd__buf_1 _11936_ (.A(_06234_),
    .X(_06240_));
 sky130_fd_sc_hd__buf_1 _11937_ (.A(_06237_),
    .X(_06241_));
 sky130_fd_sc_hd__a22o_1 _11938_ (.A1(\r1.regblock[23][25] ),
    .A2(_06240_),
    .B1(_04255_),
    .B2(_06241_),
    .X(_02422_));
 sky130_fd_sc_hd__clkbuf_1 _11939_ (.A(_06239_),
    .X(_01396_));
 sky130_fd_sc_hd__a22o_1 _11940_ (.A1(\r1.regblock[23][24] ),
    .A2(_06240_),
    .B1(_04258_),
    .B2(_06241_),
    .X(_02421_));
 sky130_fd_sc_hd__clkbuf_1 _11941_ (.A(_06239_),
    .X(_01395_));
 sky130_fd_sc_hd__a22o_1 _11942_ (.A1(\r1.regblock[23][23] ),
    .A2(_06240_),
    .B1(_04261_),
    .B2(_06241_),
    .X(_02420_));
 sky130_fd_sc_hd__buf_2 _11943_ (.A(_03909_),
    .X(_06242_));
 sky130_fd_sc_hd__buf_1 _11944_ (.A(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_1 _11945_ (.A(_06243_),
    .X(_01394_));
 sky130_fd_sc_hd__buf_1 _11946_ (.A(_06234_),
    .X(_06244_));
 sky130_fd_sc_hd__buf_1 _11947_ (.A(_06237_),
    .X(_06245_));
 sky130_fd_sc_hd__a22o_1 _11948_ (.A1(\r1.regblock[23][22] ),
    .A2(_06244_),
    .B1(_04264_),
    .B2(_06245_),
    .X(_02419_));
 sky130_fd_sc_hd__clkbuf_1 _11949_ (.A(_06243_),
    .X(_01393_));
 sky130_fd_sc_hd__a22o_1 _11950_ (.A1(\r1.regblock[23][21] ),
    .A2(_06244_),
    .B1(_04267_),
    .B2(_06245_),
    .X(_02418_));
 sky130_fd_sc_hd__clkbuf_1 _11951_ (.A(_06243_),
    .X(_01392_));
 sky130_fd_sc_hd__a22o_1 _11952_ (.A1(\r1.regblock[23][20] ),
    .A2(_06244_),
    .B1(_04271_),
    .B2(_06245_),
    .X(_02417_));
 sky130_fd_sc_hd__buf_1 _11953_ (.A(_06242_),
    .X(_06246_));
 sky130_fd_sc_hd__clkbuf_1 _11954_ (.A(_06246_),
    .X(_01391_));
 sky130_fd_sc_hd__buf_2 _11955_ (.A(_06233_),
    .X(_06247_));
 sky130_fd_sc_hd__buf_1 _11956_ (.A(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__clkbuf_2 _11957_ (.A(_06236_),
    .X(_06249_));
 sky130_fd_sc_hd__buf_1 _11958_ (.A(_06249_),
    .X(_06250_));
 sky130_fd_sc_hd__a22o_1 _11959_ (.A1(\r1.regblock[23][19] ),
    .A2(_06248_),
    .B1(_04275_),
    .B2(_06250_),
    .X(_02416_));
 sky130_fd_sc_hd__clkbuf_1 _11960_ (.A(_06246_),
    .X(_01390_));
 sky130_fd_sc_hd__a22o_1 _11961_ (.A1(\r1.regblock[23][18] ),
    .A2(_06248_),
    .B1(_04279_),
    .B2(_06250_),
    .X(_02415_));
 sky130_fd_sc_hd__clkbuf_1 _11962_ (.A(_06246_),
    .X(_01389_));
 sky130_fd_sc_hd__a22o_1 _11963_ (.A1(\r1.regblock[23][17] ),
    .A2(_06248_),
    .B1(_04282_),
    .B2(_06250_),
    .X(_02414_));
 sky130_fd_sc_hd__buf_1 _11964_ (.A(_06242_),
    .X(_06251_));
 sky130_fd_sc_hd__clkbuf_1 _11965_ (.A(_06251_),
    .X(_01388_));
 sky130_fd_sc_hd__buf_1 _11966_ (.A(_06247_),
    .X(_06252_));
 sky130_fd_sc_hd__buf_1 _11967_ (.A(_06249_),
    .X(_06253_));
 sky130_fd_sc_hd__a22o_1 _11968_ (.A1(\r1.regblock[23][16] ),
    .A2(_06252_),
    .B1(_04285_),
    .B2(_06253_),
    .X(_02413_));
 sky130_fd_sc_hd__clkbuf_1 _11969_ (.A(_06251_),
    .X(_01387_));
 sky130_fd_sc_hd__a22o_1 _11970_ (.A1(\r1.regblock[23][15] ),
    .A2(_06252_),
    .B1(_04288_),
    .B2(_06253_),
    .X(_02412_));
 sky130_fd_sc_hd__clkbuf_1 _11971_ (.A(_06251_),
    .X(_01386_));
 sky130_fd_sc_hd__a22o_1 _11972_ (.A1(\r1.regblock[23][14] ),
    .A2(_06252_),
    .B1(_04291_),
    .B2(_06253_),
    .X(_02411_));
 sky130_fd_sc_hd__clkbuf_4 _11973_ (.A(_03909_),
    .X(_06254_));
 sky130_fd_sc_hd__buf_1 _11974_ (.A(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__clkbuf_1 _11975_ (.A(_06255_),
    .X(_01385_));
 sky130_fd_sc_hd__buf_1 _11976_ (.A(_06247_),
    .X(_06256_));
 sky130_fd_sc_hd__buf_1 _11977_ (.A(_06249_),
    .X(_06257_));
 sky130_fd_sc_hd__a22o_1 _11978_ (.A1(\r1.regblock[23][13] ),
    .A2(_06256_),
    .B1(_04294_),
    .B2(_06257_),
    .X(_02410_));
 sky130_fd_sc_hd__clkbuf_1 _11979_ (.A(_06255_),
    .X(_01384_));
 sky130_fd_sc_hd__a22o_1 _11980_ (.A1(\r1.regblock[23][12] ),
    .A2(_06256_),
    .B1(_04297_),
    .B2(_06257_),
    .X(_02409_));
 sky130_fd_sc_hd__clkbuf_1 _11981_ (.A(_06255_),
    .X(_01383_));
 sky130_fd_sc_hd__a22o_1 _11982_ (.A1(\r1.regblock[23][11] ),
    .A2(_06256_),
    .B1(_04301_),
    .B2(_06257_),
    .X(_02408_));
 sky130_fd_sc_hd__buf_1 _11983_ (.A(_06254_),
    .X(_06258_));
 sky130_fd_sc_hd__clkbuf_1 _11984_ (.A(_06258_),
    .X(_01382_));
 sky130_fd_sc_hd__clkbuf_2 _11985_ (.A(_06233_),
    .X(_06259_));
 sky130_fd_sc_hd__buf_1 _11986_ (.A(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__clkbuf_2 _11987_ (.A(_06236_),
    .X(_06261_));
 sky130_fd_sc_hd__buf_1 _11988_ (.A(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__a22o_1 _11989_ (.A1(\r1.regblock[23][10] ),
    .A2(_06260_),
    .B1(_04305_),
    .B2(_06262_),
    .X(_02407_));
 sky130_fd_sc_hd__clkbuf_1 _11990_ (.A(_06258_),
    .X(_01381_));
 sky130_fd_sc_hd__a22o_1 _11991_ (.A1(\r1.regblock[23][9] ),
    .A2(_06260_),
    .B1(_04309_),
    .B2(_06262_),
    .X(_02406_));
 sky130_fd_sc_hd__clkbuf_1 _11992_ (.A(_06258_),
    .X(_01380_));
 sky130_fd_sc_hd__a22o_1 _11993_ (.A1(\r1.regblock[23][8] ),
    .A2(_06260_),
    .B1(_04312_),
    .B2(_06262_),
    .X(_02405_));
 sky130_fd_sc_hd__buf_1 _11994_ (.A(_06254_),
    .X(_06263_));
 sky130_fd_sc_hd__clkbuf_1 _11995_ (.A(_06263_),
    .X(_01379_));
 sky130_fd_sc_hd__buf_1 _11996_ (.A(_06259_),
    .X(_06264_));
 sky130_fd_sc_hd__buf_1 _11997_ (.A(_06261_),
    .X(_06265_));
 sky130_fd_sc_hd__a22o_1 _11998_ (.A1(\r1.regblock[23][7] ),
    .A2(_06264_),
    .B1(_04315_),
    .B2(_06265_),
    .X(_02404_));
 sky130_fd_sc_hd__clkbuf_1 _11999_ (.A(_06263_),
    .X(_01378_));
 sky130_fd_sc_hd__a22o_1 _12000_ (.A1(\r1.regblock[23][6] ),
    .A2(_06264_),
    .B1(_04318_),
    .B2(_06265_),
    .X(_02403_));
 sky130_fd_sc_hd__clkbuf_1 _12001_ (.A(_06263_),
    .X(_01377_));
 sky130_fd_sc_hd__a22o_1 _12002_ (.A1(\r1.regblock[23][5] ),
    .A2(_06264_),
    .B1(_04321_),
    .B2(_06265_),
    .X(_02402_));
 sky130_fd_sc_hd__buf_1 _12003_ (.A(_03910_),
    .X(_06266_));
 sky130_fd_sc_hd__clkbuf_1 _12004_ (.A(_06266_),
    .X(_01376_));
 sky130_fd_sc_hd__buf_1 _12005_ (.A(_06259_),
    .X(_06267_));
 sky130_fd_sc_hd__buf_1 _12006_ (.A(_06261_),
    .X(_06268_));
 sky130_fd_sc_hd__a22o_1 _12007_ (.A1(\r1.regblock[23][4] ),
    .A2(_06267_),
    .B1(_04324_),
    .B2(_06268_),
    .X(_02401_));
 sky130_fd_sc_hd__clkbuf_1 _12008_ (.A(_06266_),
    .X(_01375_));
 sky130_fd_sc_hd__a22o_1 _12009_ (.A1(\r1.regblock[23][3] ),
    .A2(_06267_),
    .B1(_04327_),
    .B2(_06268_),
    .X(_02400_));
 sky130_fd_sc_hd__clkbuf_1 _12010_ (.A(_06266_),
    .X(_01374_));
 sky130_fd_sc_hd__a22o_1 _12011_ (.A1(\r1.regblock[23][2] ),
    .A2(_06267_),
    .B1(_04332_),
    .B2(_06268_),
    .X(_02399_));
 sky130_fd_sc_hd__buf_1 _12012_ (.A(_03910_),
    .X(_06269_));
 sky130_fd_sc_hd__clkbuf_1 _12013_ (.A(_06269_),
    .X(_01373_));
 sky130_fd_sc_hd__a22o_1 _12014_ (.A1(\r1.regblock[23][1] ),
    .A2(_06227_),
    .B1(_04334_),
    .B2(_06230_),
    .X(_02398_));
 sky130_fd_sc_hd__clkbuf_1 _12015_ (.A(_06269_),
    .X(_01372_));
 sky130_fd_sc_hd__a22o_1 _12016_ (.A1(\r1.regblock[23][0] ),
    .A2(_06227_),
    .B1(_04336_),
    .B2(_06230_),
    .X(_02397_));
 sky130_fd_sc_hd__clkbuf_1 _12017_ (.A(_06269_),
    .X(_01371_));
 sky130_fd_sc_hd__clkbuf_1 _12018_ (.A(_03911_),
    .X(_01370_));
 sky130_fd_sc_hd__clkbuf_1 _12019_ (.A(_03911_),
    .X(_01369_));
 sky130_fd_sc_hd__buf_1 _12020_ (.A(\e1.alu1.a[24] ),
    .X(_06270_));
 sky130_fd_sc_hd__buf_1 _12021_ (.A(\e1.alu1.a1.b[24] ),
    .X(_06271_));
 sky130_fd_sc_hd__inv_2 _12022_ (.A(\c1.instruction2[4] ),
    .Y(_06272_));
 sky130_fd_sc_hd__or4_4 _12023_ (.A(\c1.instruction2[6] ),
    .B(_06272_),
    .C(\c1.instruction2[5] ),
    .D(_03678_),
    .X(_06273_));
 sky130_fd_sc_hd__buf_1 _12024_ (.A(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__or2_1 _12025_ (.A(\c1.instruction2[14] ),
    .B(_03967_),
    .X(_06275_));
 sky130_fd_sc_hd__buf_1 _12026_ (.A(_06275_),
    .X(_00005_));
 sky130_fd_sc_hd__inv_2 _12027_ (.A(_00005_),
    .Y(_06276_));
 sky130_fd_sc_hd__a31o_1 _12028_ (.A1(_03968_),
    .A2(\c1.instruction2[12] ),
    .A3(_03965_),
    .B1(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__inv_2 _12029_ (.A(_06277_),
    .Y(_00006_));
 sky130_fd_sc_hd__or4_4 _12030_ (.A(_03675_),
    .B(_06272_),
    .C(_03677_),
    .D(_03679_),
    .X(_06278_));
 sky130_fd_sc_hd__buf_1 _12031_ (.A(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__o22a_2 _12032_ (.A1(_06274_),
    .A2(_00006_),
    .B1(_00019_),
    .B2(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__inv_2 _12033_ (.A(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__clkbuf_1 _12034_ (.A(\c1.instruction2[13] ),
    .X(_06282_));
 sky130_fd_sc_hd__or2_2 _12035_ (.A(_06282_),
    .B(_03970_),
    .X(_06283_));
 sky130_fd_sc_hd__or2_2 _12036_ (.A(_03966_),
    .B(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__or2_1 _12037_ (.A(_06272_),
    .B(\c1.instruction2[29] ),
    .X(_06285_));
 sky130_fd_sc_hd__or3_1 _12038_ (.A(\c1.instruction2[28] ),
    .B(\c1.instruction2[27] ),
    .C(\c1.instruction2[31] ),
    .X(_06286_));
 sky130_fd_sc_hd__or3_4 _12039_ (.A(\c1.instruction2[26] ),
    .B(\c1.instruction2[25] ),
    .C(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__or2_2 _12040_ (.A(_03675_),
    .B(_03679_),
    .X(_06288_));
 sky130_fd_sc_hd__o21a_1 _12041_ (.A1(_03974_),
    .A2(_06288_),
    .B1(_03680_),
    .X(_06289_));
 sky130_fd_sc_hd__o41a_4 _12042_ (.A1(_06284_),
    .A2(_06285_),
    .A3(_06287_),
    .A4(_06288_),
    .B1(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__inv_2 _12043_ (.A(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__or2_1 _12044_ (.A(_06281_),
    .B(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__inv_2 _12045_ (.A(_00018_),
    .Y(_06293_));
 sky130_fd_sc_hd__o221a_2 _12046_ (.A1(_06293_),
    .A2(_06279_),
    .B1(_00015_),
    .B2(_06274_),
    .C1(_06289_),
    .X(_06294_));
 sky130_fd_sc_hd__inv_2 _12047_ (.A(_06294_),
    .Y(_06295_));
 sky130_fd_sc_hd__inv_2 _12048_ (.A(_00013_),
    .Y(_06296_));
 sky130_fd_sc_hd__buf_1 _12049_ (.A(_03964_),
    .X(_06297_));
 sky130_fd_sc_hd__nor2_4 _12050_ (.A(_06297_),
    .B(_06277_),
    .Y(_00007_));
 sky130_fd_sc_hd__or3b_2 _12051_ (.A(\c1.instruction2[29] ),
    .B(_06287_),
    .C_N(\c1.instruction2[30] ),
    .X(_06298_));
 sky130_fd_sc_hd__buf_1 _12052_ (.A(_06298_),
    .X(_00010_));
 sky130_fd_sc_hd__buf_1 _12053_ (.A(\c1.instruction2[12] ),
    .X(_06299_));
 sky130_fd_sc_hd__o21a_1 _12054_ (.A1(_03968_),
    .A2(_06299_),
    .B1(_06283_),
    .X(_06300_));
 sky130_fd_sc_hd__a31oi_2 _12055_ (.A1(_03964_),
    .A2(_03969_),
    .A3(_00010_),
    .B1(_06300_),
    .Y(_00011_));
 sky130_fd_sc_hd__o21bai_1 _12056_ (.A1(_00007_),
    .A2(_00011_),
    .B1_N(_06274_),
    .Y(_06301_));
 sky130_fd_sc_hd__o221a_2 _12057_ (.A1(_03974_),
    .A2(_06288_),
    .B1(_06296_),
    .B2(_06279_),
    .C1(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__or2_1 _12058_ (.A(_06295_),
    .B(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__or2_2 _12059_ (.A(_06292_),
    .B(_06303_),
    .X(_06304_));
 sky130_fd_sc_hd__inv_2 _12060_ (.A(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__buf_1 _12061_ (.A(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__buf_1 _12062_ (.A(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__o21a_1 _12063_ (.A1(_06270_),
    .A2(_06271_),
    .B1(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__inv_2 _12064_ (.A(\e1.alu1.a[22] ),
    .Y(_06309_));
 sky130_fd_sc_hd__buf_1 _12065_ (.A(\e1.alu1.a1.b[22] ),
    .X(_06310_));
 sky130_fd_sc_hd__o22a_1 _12066_ (.A1(_06273_),
    .A2(_00005_),
    .B1(_00098_),
    .B2(_06278_),
    .X(_06311_));
 sky130_fd_sc_hd__buf_1 _12067_ (.A(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__buf_1 _12068_ (.A(_06312_),
    .X(_06313_));
 sky130_fd_sc_hd__buf_1 _12069_ (.A(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__inv_2 _12070_ (.A(\e1.alu1.a1.b[22] ),
    .Y(_06315_));
 sky130_fd_sc_hd__inv_2 _12071_ (.A(_06311_),
    .Y(_06316_));
 sky130_fd_sc_hd__buf_1 _12072_ (.A(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__buf_1 _12073_ (.A(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__o22a_1 _12074_ (.A1(_06310_),
    .A2(_06314_),
    .B1(_06315_),
    .B2(_06318_),
    .X(_06319_));
 sky130_fd_sc_hd__or2_1 _12075_ (.A(_06309_),
    .B(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__inv_2 _12076_ (.A(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__a21oi_2 _12077_ (.A1(_06309_),
    .A2(_06319_),
    .B1(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__clkbuf_2 _12078_ (.A(\e1.alu1.a[23] ),
    .X(_06323_));
 sky130_fd_sc_hd__buf_1 _12079_ (.A(\e1.alu1.a1.b[23] ),
    .X(_06324_));
 sky130_fd_sc_hd__buf_1 _12080_ (.A(_06312_),
    .X(_06325_));
 sky130_fd_sc_hd__buf_1 _12081_ (.A(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__clkbuf_2 _12082_ (.A(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__inv_2 _12083_ (.A(\e1.alu1.a1.b[23] ),
    .Y(_06328_));
 sky130_fd_sc_hd__clkbuf_2 _12084_ (.A(_06318_),
    .X(_06329_));
 sky130_fd_sc_hd__o22a_1 _12085_ (.A1(_06324_),
    .A2(_06327_),
    .B1(_06328_),
    .B2(_06329_),
    .X(_06330_));
 sky130_fd_sc_hd__inv_2 _12086_ (.A(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__nor2_2 _12087_ (.A(\e1.alu1.a[23] ),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__a21oi_4 _12088_ (.A1(_06323_),
    .A2(_06331_),
    .B1(_06332_),
    .Y(_06333_));
 sky130_fd_sc_hd__nand2_1 _12089_ (.A(_06322_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__inv_2 _12090_ (.A(\e1.alu1.a[20] ),
    .Y(_06335_));
 sky130_fd_sc_hd__buf_1 _12091_ (.A(\e1.alu1.a1.b[20] ),
    .X(_06336_));
 sky130_fd_sc_hd__buf_1 _12092_ (.A(_06314_),
    .X(_06337_));
 sky130_fd_sc_hd__inv_2 _12093_ (.A(\e1.alu1.a1.b[20] ),
    .Y(_06338_));
 sky130_fd_sc_hd__clkbuf_2 _12094_ (.A(_06318_),
    .X(_06339_));
 sky130_fd_sc_hd__o22a_1 _12095_ (.A1(_06336_),
    .A2(_06337_),
    .B1(_06338_),
    .B2(_06339_),
    .X(_06340_));
 sky130_fd_sc_hd__buf_1 _12096_ (.A(\e1.alu1.a[20] ),
    .X(_06341_));
 sky130_fd_sc_hd__inv_2 _12097_ (.A(_06340_),
    .Y(_06342_));
 sky130_fd_sc_hd__o22a_1 _12098_ (.A1(_06335_),
    .A2(_06340_),
    .B1(_06341_),
    .B2(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__inv_2 _12099_ (.A(\e1.alu1.a[21] ),
    .Y(_06344_));
 sky130_fd_sc_hd__buf_1 _12100_ (.A(_06344_),
    .X(_06345_));
 sky130_fd_sc_hd__buf_1 _12101_ (.A(\e1.alu1.a1.b[21] ),
    .X(_06346_));
 sky130_fd_sc_hd__buf_1 _12102_ (.A(_06326_),
    .X(_06347_));
 sky130_fd_sc_hd__buf_1 _12103_ (.A(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__inv_2 _12104_ (.A(\e1.alu1.a1.b[21] ),
    .Y(_06349_));
 sky130_fd_sc_hd__buf_1 _12105_ (.A(_06317_),
    .X(_06350_));
 sky130_fd_sc_hd__buf_1 _12106_ (.A(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__buf_1 _12107_ (.A(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__o22a_1 _12108_ (.A1(_06346_),
    .A2(_06348_),
    .B1(_06349_),
    .B2(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__nor2_1 _12109_ (.A(_06344_),
    .B(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__a21oi_2 _12110_ (.A1(_06345_),
    .A2(_06353_),
    .B1(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__nand3b_2 _12111_ (.A_N(_06334_),
    .B(_06343_),
    .C(_06355_),
    .Y(_06356_));
 sky130_fd_sc_hd__inv_2 _12112_ (.A(\e1.alu1.a[19] ),
    .Y(_06357_));
 sky130_fd_sc_hd__buf_1 _12113_ (.A(\e1.alu1.a1.b[19] ),
    .X(_06358_));
 sky130_fd_sc_hd__inv_2 _12114_ (.A(\e1.alu1.a1.b[19] ),
    .Y(_06359_));
 sky130_fd_sc_hd__o22a_1 _12115_ (.A1(_06358_),
    .A2(_06347_),
    .B1(_06359_),
    .B2(_06329_),
    .X(_06360_));
 sky130_fd_sc_hd__buf_1 _12116_ (.A(\e1.alu1.a[19] ),
    .X(_06361_));
 sky130_fd_sc_hd__inv_2 _12117_ (.A(_06360_),
    .Y(_06362_));
 sky130_fd_sc_hd__o22a_1 _12118_ (.A1(_06357_),
    .A2(_06360_),
    .B1(_06361_),
    .B2(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__inv_2 _12119_ (.A(\e1.alu1.a[18] ),
    .Y(_06364_));
 sky130_fd_sc_hd__buf_1 _12120_ (.A(\e1.alu1.a1.b[18] ),
    .X(_06365_));
 sky130_fd_sc_hd__inv_2 _12121_ (.A(\e1.alu1.a1.b[18] ),
    .Y(_06366_));
 sky130_fd_sc_hd__o22a_1 _12122_ (.A1(_06365_),
    .A2(_06337_),
    .B1(_06366_),
    .B2(_06352_),
    .X(_06367_));
 sky130_fd_sc_hd__nor2_1 _12123_ (.A(_06364_),
    .B(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__a21oi_2 _12124_ (.A1(_06364_),
    .A2(_06367_),
    .B1(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__nand2_1 _12125_ (.A(_06363_),
    .B(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__inv_2 _12126_ (.A(\e1.alu1.a[16] ),
    .Y(_06371_));
 sky130_fd_sc_hd__inv_2 _12127_ (.A(\e1.alu1.a1.b[16] ),
    .Y(_06372_));
 sky130_fd_sc_hd__buf_1 _12128_ (.A(_06316_),
    .X(_06373_));
 sky130_fd_sc_hd__buf_1 _12129_ (.A(_06373_),
    .X(_06374_));
 sky130_fd_sc_hd__clkbuf_2 _12130_ (.A(_06374_),
    .X(_06375_));
 sky130_fd_sc_hd__o22a_1 _12131_ (.A1(\e1.alu1.a1.b[16] ),
    .A2(_06314_),
    .B1(_06372_),
    .B2(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__buf_1 _12132_ (.A(\e1.alu1.a[16] ),
    .X(_06377_));
 sky130_fd_sc_hd__inv_2 _12133_ (.A(_06376_),
    .Y(_06378_));
 sky130_fd_sc_hd__o22a_1 _12134_ (.A1(_06371_),
    .A2(_06376_),
    .B1(_06377_),
    .B2(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__inv_2 _12135_ (.A(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__inv_2 _12136_ (.A(\e1.alu1.a[17] ),
    .Y(_06381_));
 sky130_fd_sc_hd__buf_1 _12137_ (.A(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__clkbuf_4 _12138_ (.A(_06382_),
    .X(_00063_));
 sky130_fd_sc_hd__buf_1 _12139_ (.A(\e1.alu1.a1.b[17] ),
    .X(_06383_));
 sky130_fd_sc_hd__inv_2 _12140_ (.A(\e1.alu1.a1.b[17] ),
    .Y(_06384_));
 sky130_fd_sc_hd__o22a_1 _12141_ (.A1(_06383_),
    .A2(_06327_),
    .B1(_06384_),
    .B2(_06351_),
    .X(_06385_));
 sky130_fd_sc_hd__nor2_1 _12142_ (.A(_06381_),
    .B(_06385_),
    .Y(_06386_));
 sky130_fd_sc_hd__a21oi_1 _12143_ (.A1(_00063_),
    .A2(_06385_),
    .B1(_06386_),
    .Y(_06387_));
 sky130_fd_sc_hd__or3b_4 _12144_ (.A(_06370_),
    .B(_06380_),
    .C_N(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__clkbuf_2 _12145_ (.A(\e1.alu1.a[15] ),
    .X(_06389_));
 sky130_fd_sc_hd__buf_1 _12146_ (.A(\e1.alu1.a1.b[15] ),
    .X(_06390_));
 sky130_fd_sc_hd__inv_2 _12147_ (.A(\e1.alu1.a1.b[15] ),
    .Y(_06391_));
 sky130_fd_sc_hd__buf_1 _12148_ (.A(_06373_),
    .X(_06392_));
 sky130_fd_sc_hd__o22a_1 _12149_ (.A1(_06390_),
    .A2(_06313_),
    .B1(_06391_),
    .B2(_06392_),
    .X(_06393_));
 sky130_fd_sc_hd__inv_2 _12150_ (.A(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__nor2_2 _12151_ (.A(\e1.alu1.a[15] ),
    .B(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__a21oi_4 _12152_ (.A1(_06389_),
    .A2(_06394_),
    .B1(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__inv_2 _12153_ (.A(\e1.alu1.a[14] ),
    .Y(_06397_));
 sky130_fd_sc_hd__buf_1 _12154_ (.A(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__clkbuf_2 _12155_ (.A(\e1.alu1.a1.b[14] ),
    .X(_06399_));
 sky130_fd_sc_hd__buf_1 _12156_ (.A(_06312_),
    .X(_06400_));
 sky130_fd_sc_hd__buf_1 _12157_ (.A(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__inv_2 _12158_ (.A(\e1.alu1.a1.b[14] ),
    .Y(_06402_));
 sky130_fd_sc_hd__o22a_1 _12159_ (.A1(_06399_),
    .A2(_06401_),
    .B1(_06402_),
    .B2(_06392_),
    .X(_06403_));
 sky130_fd_sc_hd__or2_1 _12160_ (.A(_06397_),
    .B(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__a21boi_4 _12161_ (.A1(_06398_),
    .A2(_06403_),
    .B1_N(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand2_1 _12162_ (.A(_06396_),
    .B(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__inv_2 _12163_ (.A(\e1.alu1.a[12] ),
    .Y(_06407_));
 sky130_fd_sc_hd__clkbuf_2 _12164_ (.A(_06313_),
    .X(_06408_));
 sky130_fd_sc_hd__inv_2 _12165_ (.A(\e1.alu1.a1.b[12] ),
    .Y(_06409_));
 sky130_fd_sc_hd__o22a_1 _12166_ (.A1(\e1.alu1.a1.b[12] ),
    .A2(_06408_),
    .B1(_06409_),
    .B2(_06375_),
    .X(_06410_));
 sky130_fd_sc_hd__buf_1 _12167_ (.A(\e1.alu1.a[12] ),
    .X(_06411_));
 sky130_fd_sc_hd__inv_2 _12168_ (.A(_06410_),
    .Y(_06412_));
 sky130_fd_sc_hd__o22a_1 _12169_ (.A1(_06407_),
    .A2(_06410_),
    .B1(_06411_),
    .B2(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__inv_2 _12170_ (.A(\e1.alu1.a[13] ),
    .Y(_06414_));
 sky130_fd_sc_hd__buf_1 _12171_ (.A(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__buf_1 _12172_ (.A(\e1.alu1.a1.b[13] ),
    .X(_06416_));
 sky130_fd_sc_hd__inv_2 _12173_ (.A(\e1.alu1.a1.b[13] ),
    .Y(_06417_));
 sky130_fd_sc_hd__o22a_1 _12174_ (.A1(_06416_),
    .A2(_06327_),
    .B1(_06417_),
    .B2(_06329_),
    .X(_06418_));
 sky130_fd_sc_hd__nor2_1 _12175_ (.A(_06414_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__a21oi_2 _12176_ (.A1(_06415_),
    .A2(_06418_),
    .B1(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__nand3b_2 _12177_ (.A_N(_06406_),
    .B(_06413_),
    .C(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__inv_2 _12178_ (.A(\e1.alu1.a[11] ),
    .Y(_06422_));
 sky130_fd_sc_hd__buf_1 _12179_ (.A(\e1.alu1.a1.b[11] ),
    .X(_06423_));
 sky130_fd_sc_hd__inv_2 _12180_ (.A(\e1.alu1.a1.b[11] ),
    .Y(_06424_));
 sky130_fd_sc_hd__o22a_1 _12181_ (.A1(_06423_),
    .A2(_06326_),
    .B1(_06424_),
    .B2(_06350_),
    .X(_06425_));
 sky130_fd_sc_hd__buf_1 _12182_ (.A(\e1.alu1.a[11] ),
    .X(_06426_));
 sky130_fd_sc_hd__inv_2 _12183_ (.A(_06425_),
    .Y(_06427_));
 sky130_fd_sc_hd__o22a_1 _12184_ (.A1(_06422_),
    .A2(_06425_),
    .B1(_06426_),
    .B2(_06427_),
    .X(_06428_));
 sky130_fd_sc_hd__inv_2 _12185_ (.A(\e1.alu1.a[10] ),
    .Y(_06429_));
 sky130_fd_sc_hd__clkbuf_2 _12186_ (.A(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__clkbuf_2 _12187_ (.A(\e1.alu1.a1.b[10] ),
    .X(_06431_));
 sky130_fd_sc_hd__inv_2 _12188_ (.A(\e1.alu1.a1.b[10] ),
    .Y(_06432_));
 sky130_fd_sc_hd__o22a_1 _12189_ (.A1(_06431_),
    .A2(_06400_),
    .B1(_06432_),
    .B2(_06373_),
    .X(_06433_));
 sky130_fd_sc_hd__or2_1 _12190_ (.A(_06429_),
    .B(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__inv_2 _12191_ (.A(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__a21oi_4 _12192_ (.A1(_06430_),
    .A2(_06433_),
    .B1(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__nand2_1 _12193_ (.A(_06428_),
    .B(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__inv_2 _12194_ (.A(\e1.alu1.a[8] ),
    .Y(_06438_));
 sky130_fd_sc_hd__clkbuf_2 _12195_ (.A(\e1.alu1.a1.b[8] ),
    .X(_06439_));
 sky130_fd_sc_hd__inv_2 _12196_ (.A(\e1.alu1.a1.b[8] ),
    .Y(_06440_));
 sky130_fd_sc_hd__o22a_1 _12197_ (.A1(_06439_),
    .A2(_06325_),
    .B1(_06440_),
    .B2(_06374_),
    .X(_06441_));
 sky130_fd_sc_hd__buf_1 _12198_ (.A(\e1.alu1.a[8] ),
    .X(_06442_));
 sky130_fd_sc_hd__inv_2 _12199_ (.A(_06441_),
    .Y(_06443_));
 sky130_fd_sc_hd__o22a_1 _12200_ (.A1(_06438_),
    .A2(_06441_),
    .B1(_06442_),
    .B2(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__inv_2 _12201_ (.A(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__inv_2 _12202_ (.A(\e1.alu1.a[9] ),
    .Y(_06446_));
 sky130_fd_sc_hd__buf_1 _12203_ (.A(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__buf_1 _12204_ (.A(\e1.alu1.a1.b[9] ),
    .X(_06448_));
 sky130_fd_sc_hd__inv_2 _12205_ (.A(\e1.alu1.a1.b[9] ),
    .Y(_06449_));
 sky130_fd_sc_hd__o22a_1 _12206_ (.A1(_06448_),
    .A2(_06401_),
    .B1(_06449_),
    .B2(_06392_),
    .X(_06450_));
 sky130_fd_sc_hd__nor2_1 _12207_ (.A(_06446_),
    .B(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__a21oi_1 _12208_ (.A1(_06447_),
    .A2(_06450_),
    .B1(_06451_),
    .Y(_06452_));
 sky130_fd_sc_hd__or3b_1 _12209_ (.A(_06437_),
    .B(_06445_),
    .C_N(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__inv_2 _12210_ (.A(\e1.alu1.a[3] ),
    .Y(_06454_));
 sky130_fd_sc_hd__clkbuf_4 _12211_ (.A(_06454_),
    .X(_00035_));
 sky130_fd_sc_hd__buf_1 _12212_ (.A(\e1.alu1.a1.b[3] ),
    .X(_06455_));
 sky130_fd_sc_hd__inv_2 _12213_ (.A(\e1.alu1.a1.b[3] ),
    .Y(_06456_));
 sky130_fd_sc_hd__o22a_2 _12214_ (.A1(_06455_),
    .A2(_06337_),
    .B1(_06456_),
    .B2(_06339_),
    .X(_06457_));
 sky130_fd_sc_hd__nor2_2 _12215_ (.A(_06454_),
    .B(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__a21oi_4 _12216_ (.A1(_00035_),
    .A2(_06457_),
    .B1(_06458_),
    .Y(_06459_));
 sky130_fd_sc_hd__inv_2 _12217_ (.A(\e1.alu1.a[2] ),
    .Y(_06460_));
 sky130_fd_sc_hd__inv_2 _12218_ (.A(\e1.alu1.a1.b[2] ),
    .Y(_06461_));
 sky130_fd_sc_hd__o22a_1 _12219_ (.A1(\e1.alu1.a1.b[2] ),
    .A2(_06408_),
    .B1(_06461_),
    .B2(_06351_),
    .X(_06462_));
 sky130_fd_sc_hd__inv_2 _12220_ (.A(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__o22a_1 _12221_ (.A1(_06460_),
    .A2(_06462_),
    .B1(\e1.alu1.a[2] ),
    .B2(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__inv_2 _12222_ (.A(\e1.alu1.a[1] ),
    .Y(_06465_));
 sky130_fd_sc_hd__buf_1 _12223_ (.A(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__inv_2 _12224_ (.A(\e1.alu1.a1.b[1] ),
    .Y(_06467_));
 sky130_fd_sc_hd__o22a_1 _12225_ (.A1(\e1.alu1.a1.b[1] ),
    .A2(_06401_),
    .B1(_06467_),
    .B2(_06350_),
    .X(_06468_));
 sky130_fd_sc_hd__a2bb2o_1 _12226_ (.A1_N(_06465_),
    .A2_N(_06468_),
    .B1(_06465_),
    .B2(_06468_),
    .X(_06469_));
 sky130_fd_sc_hd__o22a_1 _12227_ (.A1(_06466_),
    .A2(_06468_),
    .B1(_00135_),
    .B2(_06469_),
    .X(_06470_));
 sky130_fd_sc_hd__inv_2 _12228_ (.A(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__buf_1 _12229_ (.A(\e1.alu1.a[2] ),
    .X(_06472_));
 sky130_fd_sc_hd__nand2_1 _12230_ (.A(_06454_),
    .B(_06457_),
    .Y(_06473_));
 sky130_fd_sc_hd__a31o_1 _12231_ (.A1(_06472_),
    .A2(_06463_),
    .A3(_06473_),
    .B1(_06458_),
    .X(_06474_));
 sky130_fd_sc_hd__a31o_1 _12232_ (.A1(_06459_),
    .A2(_06464_),
    .A3(_06471_),
    .B1(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__buf_1 _12233_ (.A(\e1.alu1.a[7] ),
    .X(_06476_));
 sky130_fd_sc_hd__inv_2 _12234_ (.A(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__buf_1 _12235_ (.A(\e1.alu1.a1.b[7] ),
    .X(_06478_));
 sky130_fd_sc_hd__inv_2 _12236_ (.A(\e1.alu1.a1.b[7] ),
    .Y(_06479_));
 sky130_fd_sc_hd__o22a_1 _12237_ (.A1(_06478_),
    .A2(_06400_),
    .B1(_06479_),
    .B2(_06317_),
    .X(_06480_));
 sky130_fd_sc_hd__inv_2 _12238_ (.A(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__or2_1 _12239_ (.A(\e1.alu1.a[7] ),
    .B(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__o21a_1 _12240_ (.A1(_06477_),
    .A2(_06480_),
    .B1(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__inv_2 _12241_ (.A(\e1.alu1.a[6] ),
    .Y(_06484_));
 sky130_fd_sc_hd__buf_1 _12242_ (.A(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__clkbuf_2 _12243_ (.A(\e1.alu1.a1.b[6] ),
    .X(_06486_));
 sky130_fd_sc_hd__inv_2 _12244_ (.A(\e1.alu1.a1.b[6] ),
    .Y(_06487_));
 sky130_fd_sc_hd__o22a_1 _12245_ (.A1(_06486_),
    .A2(_06325_),
    .B1(_06487_),
    .B2(_06374_),
    .X(_06488_));
 sky130_fd_sc_hd__or2_1 _12246_ (.A(_06484_),
    .B(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__inv_2 _12247_ (.A(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__a21oi_1 _12248_ (.A1(_06485_),
    .A2(_06488_),
    .B1(_06490_),
    .Y(_06491_));
 sky130_fd_sc_hd__inv_2 _12249_ (.A(\e1.alu1.a[5] ),
    .Y(_06492_));
 sky130_fd_sc_hd__buf_1 _12250_ (.A(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__buf_1 _12251_ (.A(\e1.alu1.a1.b[5] ),
    .X(_06494_));
 sky130_fd_sc_hd__inv_2 _12252_ (.A(\e1.alu1.a1.b[5] ),
    .Y(_06495_));
 sky130_fd_sc_hd__o22a_1 _12253_ (.A1(_06494_),
    .A2(_06347_),
    .B1(_06495_),
    .B2(_06339_),
    .X(_06496_));
 sky130_fd_sc_hd__nor2_1 _12254_ (.A(_06492_),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__a21oi_1 _12255_ (.A1(_06493_),
    .A2(_06496_),
    .B1(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__inv_2 _12256_ (.A(\e1.alu1.a[4] ),
    .Y(_06499_));
 sky130_fd_sc_hd__buf_1 _12257_ (.A(\e1.alu1.a1.b[4] ),
    .X(_06500_));
 sky130_fd_sc_hd__inv_2 _12258_ (.A(\e1.alu1.a1.b[4] ),
    .Y(_06501_));
 sky130_fd_sc_hd__o22a_1 _12259_ (.A1(_06500_),
    .A2(_06408_),
    .B1(_06501_),
    .B2(_06375_),
    .X(_06502_));
 sky130_fd_sc_hd__buf_1 _12260_ (.A(\e1.alu1.a[4] ),
    .X(_06503_));
 sky130_fd_sc_hd__inv_2 _12261_ (.A(_06502_),
    .Y(_06504_));
 sky130_fd_sc_hd__o22a_1 _12262_ (.A1(_06499_),
    .A2(_06502_),
    .B1(_06503_),
    .B2(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__and4_1 _12263_ (.A(_06483_),
    .B(_06491_),
    .C(_06498_),
    .D(_06505_),
    .X(_06506_));
 sky130_fd_sc_hd__buf_1 _12264_ (.A(_06483_),
    .X(_06507_));
 sky130_fd_sc_hd__clkbuf_2 _12265_ (.A(_06491_),
    .X(_06508_));
 sky130_fd_sc_hd__nand2_1 _12266_ (.A(_06493_),
    .B(_06496_),
    .Y(_06509_));
 sky130_fd_sc_hd__a31o_1 _12267_ (.A1(_06503_),
    .A2(_06504_),
    .A3(_06509_),
    .B1(_06497_),
    .X(_06510_));
 sky130_fd_sc_hd__a22o_1 _12268_ (.A1(_06476_),
    .A2(_06481_),
    .B1(_06482_),
    .B2(_06490_),
    .X(_06511_));
 sky130_fd_sc_hd__a31o_1 _12269_ (.A1(_06507_),
    .A2(_06508_),
    .A3(_06510_),
    .B1(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__a21oi_4 _12270_ (.A1(_06475_),
    .A2(_06506_),
    .B1(_06512_),
    .Y(_06513_));
 sky130_fd_sc_hd__nand2_1 _12271_ (.A(_06414_),
    .B(_06418_),
    .Y(_06514_));
 sky130_fd_sc_hd__a31o_1 _12272_ (.A1(\e1.alu1.a[12] ),
    .A2(_06412_),
    .A3(_06514_),
    .B1(_06419_),
    .X(_06515_));
 sky130_fd_sc_hd__inv_2 _12273_ (.A(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__buf_1 _12274_ (.A(_06422_),
    .X(_06517_));
 sky130_fd_sc_hd__nand2_1 _12275_ (.A(_06446_),
    .B(_06450_),
    .Y(_06518_));
 sky130_fd_sc_hd__a31o_1 _12276_ (.A1(_06442_),
    .A2(_06443_),
    .A3(_06518_),
    .B1(_06451_),
    .X(_06519_));
 sky130_fd_sc_hd__inv_2 _12277_ (.A(_06519_),
    .Y(_06520_));
 sky130_fd_sc_hd__o21ai_1 _12278_ (.A1(_06426_),
    .A2(_06427_),
    .B1(_06435_),
    .Y(_06521_));
 sky130_fd_sc_hd__o221a_1 _12279_ (.A1(_06517_),
    .A2(_06425_),
    .B1(_06437_),
    .B2(_06520_),
    .C1(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__inv_2 _12280_ (.A(_06389_),
    .Y(_06523_));
 sky130_fd_sc_hd__o22a_1 _12281_ (.A1(_06523_),
    .A2(_06393_),
    .B1(_06395_),
    .B2(_06404_),
    .X(_06524_));
 sky130_fd_sc_hd__o221a_1 _12282_ (.A1(_06406_),
    .A2(_06516_),
    .B1(_06421_),
    .B2(_06522_),
    .C1(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__o31a_2 _12283_ (.A1(_06421_),
    .A2(_06453_),
    .A3(_06513_),
    .B1(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__nand2_1 _12284_ (.A(_06345_),
    .B(_06353_),
    .Y(_06527_));
 sky130_fd_sc_hd__a31o_1 _12285_ (.A1(_06341_),
    .A2(_06342_),
    .A3(_06527_),
    .B1(_06354_),
    .X(_06528_));
 sky130_fd_sc_hd__inv_2 _12286_ (.A(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__nand2_1 _12287_ (.A(_06382_),
    .B(_06385_),
    .Y(_06530_));
 sky130_fd_sc_hd__a31o_1 _12288_ (.A1(\e1.alu1.a[16] ),
    .A2(_06378_),
    .A3(_06530_),
    .B1(_06386_),
    .X(_06531_));
 sky130_fd_sc_hd__inv_2 _12289_ (.A(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__buf_1 _12290_ (.A(_06368_),
    .X(_06533_));
 sky130_fd_sc_hd__o21ai_1 _12291_ (.A1(_06361_),
    .A2(_06362_),
    .B1(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__o221a_1 _12292_ (.A1(_06357_),
    .A2(_06360_),
    .B1(_06370_),
    .B2(_06532_),
    .C1(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__inv_2 _12293_ (.A(_06323_),
    .Y(_06536_));
 sky130_fd_sc_hd__o22a_1 _12294_ (.A1(_06536_),
    .A2(_06330_),
    .B1(_06320_),
    .B2(_06332_),
    .X(_06537_));
 sky130_fd_sc_hd__o221a_1 _12295_ (.A1(_06334_),
    .A2(_06529_),
    .B1(_06356_),
    .B2(_06535_),
    .C1(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__o31a_2 _12296_ (.A1(_06356_),
    .A2(_06388_),
    .A3(_06526_),
    .B1(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__inv_2 _12297_ (.A(\e1.alu1.a[24] ),
    .Y(_06540_));
 sky130_fd_sc_hd__buf_1 _12298_ (.A(_06348_),
    .X(_06541_));
 sky130_fd_sc_hd__inv_2 _12299_ (.A(\e1.alu1.a1.b[24] ),
    .Y(_06542_));
 sky130_fd_sc_hd__buf_1 _12300_ (.A(_06352_),
    .X(_06543_));
 sky130_fd_sc_hd__buf_1 _12301_ (.A(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__o22a_1 _12302_ (.A1(_06271_),
    .A2(_06541_),
    .B1(_06542_),
    .B2(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__nor2_4 _12303_ (.A(_06540_),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__a21o_1 _12304_ (.A1(_06540_),
    .A2(_06545_),
    .B1(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__inv_2 _12305_ (.A(_06302_),
    .Y(_06548_));
 sky130_fd_sc_hd__or2_1 _12306_ (.A(_06295_),
    .B(_06548_),
    .X(_06549_));
 sky130_fd_sc_hd__or2_1 _12307_ (.A(_06294_),
    .B(_06302_),
    .X(_06550_));
 sky130_fd_sc_hd__and2_2 _12308_ (.A(_06280_),
    .B(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__a211o_1 _12309_ (.A1(_06281_),
    .A2(_06549_),
    .B1(_06291_),
    .C1(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__buf_1 _12310_ (.A(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__buf_1 _12311_ (.A(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__buf_2 _12312_ (.A(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__nor2_2 _12313_ (.A(_06539_),
    .B(_06547_),
    .Y(_06556_));
 sky130_fd_sc_hd__a211oi_4 _12314_ (.A1(_06539_),
    .A2(_06547_),
    .B1(_06555_),
    .C1(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__buf_1 _12315_ (.A(_06500_),
    .X(_06558_));
 sky130_fd_sc_hd__or3_4 _12316_ (.A(_06281_),
    .B(_06295_),
    .C(_06290_),
    .X(_06559_));
 sky130_fd_sc_hd__or2_1 _12317_ (.A(_06558_),
    .B(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__clkbuf_1 _12318_ (.A(_06560_),
    .X(_06561_));
 sky130_fd_sc_hd__buf_1 _12319_ (.A(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__buf_1 _12320_ (.A(_06455_),
    .X(_06563_));
 sky130_fd_sc_hd__buf_1 _12321_ (.A(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__clkbuf_1 _12322_ (.A(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__or2_2 _12323_ (.A(_06565_),
    .B(_00091_),
    .X(_00228_));
 sky130_fd_sc_hd__or2_1 _12324_ (.A(_06294_),
    .B(_06548_),
    .X(_06566_));
 sky130_fd_sc_hd__or2_1 _12325_ (.A(_06292_),
    .B(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__inv_2 _12326_ (.A(_06567_),
    .Y(_06568_));
 sky130_fd_sc_hd__buf_1 _12327_ (.A(_06568_),
    .X(_06569_));
 sky130_fd_sc_hd__clkbuf_2 _12328_ (.A(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__buf_4 _12329_ (.A(_06540_),
    .X(_00077_));
 sky130_fd_sc_hd__buf_1 _12330_ (.A(_06542_),
    .X(_06571_));
 sky130_fd_sc_hd__o22a_1 _12331_ (.A1(_06270_),
    .A2(_06271_),
    .B1(_00077_),
    .B2(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__a2bb2o_1 _12332_ (.A1_N(_06562_),
    .A2_N(_00228_),
    .B1(_06570_),
    .B2(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__or2_2 _12333_ (.A(_06549_),
    .B(_06292_),
    .X(_06574_));
 sky130_fd_sc_hd__buf_1 _12334_ (.A(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__buf_1 _12335_ (.A(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__buf_1 _12336_ (.A(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__or2_1 _12337_ (.A(_06280_),
    .B(_06291_),
    .X(_06578_));
 sky130_fd_sc_hd__or2_2 _12338_ (.A(_06550_),
    .B(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__buf_1 _12339_ (.A(_06579_),
    .X(_06580_));
 sky130_fd_sc_hd__buf_1 _12340_ (.A(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__o32a_1 _12341_ (.A1(_00077_),
    .A2(_06571_),
    .A3(_06577_),
    .B1(_00350_),
    .B2(_06581_),
    .X(_06582_));
 sky130_fd_sc_hd__or4b_4 _12342_ (.A(_06308_),
    .B(_06557_),
    .C(_06573_),
    .D_N(_06582_),
    .X(_00351_));
 sky130_fd_sc_hd__buf_1 _12343_ (.A(_06563_),
    .X(_06583_));
 sky130_fd_sc_hd__buf_1 _12344_ (.A(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__or2_2 _12345_ (.A(_06584_),
    .B(_00128_),
    .X(_00237_));
 sky130_fd_sc_hd__buf_1 _12346_ (.A(_06348_),
    .X(_06585_));
 sky130_fd_sc_hd__buf_1 _12347_ (.A(_06585_),
    .X(_00134_));
 sky130_fd_sc_hd__buf_1 _12348_ (.A(_06554_),
    .X(_06586_));
 sky130_fd_sc_hd__clkbuf_4 _12349_ (.A(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__inv_2 _12350_ (.A(\e1.alu1.a[25] ),
    .Y(_06588_));
 sky130_fd_sc_hd__buf_1 _12351_ (.A(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__buf_1 _12352_ (.A(\e1.alu1.a1.b[25] ),
    .X(_06590_));
 sky130_fd_sc_hd__inv_2 _12353_ (.A(\e1.alu1.a1.b[25] ),
    .Y(_06591_));
 sky130_fd_sc_hd__o22a_2 _12354_ (.A1(_06590_),
    .A2(_06541_),
    .B1(_06591_),
    .B2(_06543_),
    .X(_06592_));
 sky130_fd_sc_hd__nor2_4 _12355_ (.A(_06588_),
    .B(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__a21o_1 _12356_ (.A1(_06589_),
    .A2(_06592_),
    .B1(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__or2_1 _12357_ (.A(_06546_),
    .B(_06556_),
    .X(_06595_));
 sky130_fd_sc_hd__o2bb2a_1 _12358_ (.A1_N(_06594_),
    .A2_N(_06595_),
    .B1(_06594_),
    .B2(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__buf_1 _12359_ (.A(\e1.alu1.a[25] ),
    .X(_06597_));
 sky130_fd_sc_hd__clkbuf_2 _12360_ (.A(_06307_),
    .X(_06598_));
 sky130_fd_sc_hd__o21ai_2 _12361_ (.A1(_06590_),
    .A2(_06597_),
    .B1(_06598_),
    .Y(_06599_));
 sky130_fd_sc_hd__buf_1 _12362_ (.A(_06591_),
    .X(_06600_));
 sky130_fd_sc_hd__buf_4 _12363_ (.A(_06589_),
    .X(_00078_));
 sky130_fd_sc_hd__buf_1 _12364_ (.A(_06574_),
    .X(_06601_));
 sky130_fd_sc_hd__clkbuf_2 _12365_ (.A(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__o32a_2 _12366_ (.A1(_06600_),
    .A2(_00078_),
    .A3(_06602_),
    .B1(_00356_),
    .B2(_06581_),
    .X(_06603_));
 sky130_fd_sc_hd__buf_1 _12367_ (.A(_06560_),
    .X(_06604_));
 sky130_fd_sc_hd__buf_1 _12368_ (.A(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__buf_1 _12369_ (.A(_06567_),
    .X(_06606_));
 sky130_fd_sc_hd__buf_1 _12370_ (.A(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__clkbuf_2 _12371_ (.A(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__o22a_1 _12372_ (.A1(_06590_),
    .A2(_06597_),
    .B1(_06600_),
    .B2(_06589_),
    .X(_06609_));
 sky130_fd_sc_hd__inv_2 _12373_ (.A(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__o22a_1 _12374_ (.A1(_06605_),
    .A2(_00237_),
    .B1(_06608_),
    .B2(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__o2111ai_4 _12375_ (.A1(_06587_),
    .A2(_06596_),
    .B1(_06599_),
    .C1(_06603_),
    .D1(_06611_),
    .Y(_00357_));
 sky130_fd_sc_hd__or2_2 _12376_ (.A(_06584_),
    .B(_00149_),
    .X(_00246_));
 sky130_fd_sc_hd__buf_1 _12377_ (.A(\e1.alu1.a1.b[26] ),
    .X(_06612_));
 sky130_fd_sc_hd__clkbuf_2 _12378_ (.A(\e1.alu1.a[26] ),
    .X(_06613_));
 sky130_fd_sc_hd__nor2_2 _12379_ (.A(_06612_),
    .B(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__a21oi_2 _12380_ (.A1(_06612_),
    .A2(_06613_),
    .B1(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__inv_2 _12381_ (.A(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__buf_1 _12382_ (.A(_06579_),
    .X(_06617_));
 sky130_fd_sc_hd__buf_1 _12383_ (.A(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__buf_1 _12384_ (.A(_06304_),
    .X(_06619_));
 sky130_fd_sc_hd__o22a_1 _12385_ (.A1(_00362_),
    .A2(_06618_),
    .B1(_06619_),
    .B2(_06614_),
    .X(_06620_));
 sky130_fd_sc_hd__inv_2 _12386_ (.A(\e1.alu1.a1.b[26] ),
    .Y(_06621_));
 sky130_fd_sc_hd__inv_2 _12387_ (.A(\e1.alu1.a[26] ),
    .Y(_06622_));
 sky130_fd_sc_hd__buf_4 _12388_ (.A(_06622_),
    .X(_00080_));
 sky130_fd_sc_hd__buf_1 _12389_ (.A(_06561_),
    .X(_06623_));
 sky130_fd_sc_hd__o32a_1 _12390_ (.A1(_06621_),
    .A2(_00080_),
    .A3(_06602_),
    .B1(_06623_),
    .B2(_00246_),
    .X(_06624_));
 sky130_fd_sc_hd__o22a_2 _12391_ (.A1(_06612_),
    .A2(_06585_),
    .B1(_06621_),
    .B2(_06544_),
    .X(_06625_));
 sky130_fd_sc_hd__nor2_2 _12392_ (.A(_06622_),
    .B(_06625_),
    .Y(_06626_));
 sky130_fd_sc_hd__a21oi_4 _12393_ (.A1(_00080_),
    .A2(_06625_),
    .B1(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__inv_2 _12394_ (.A(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__nand2_2 _12395_ (.A(_00078_),
    .B(_06592_),
    .Y(_06629_));
 sky130_fd_sc_hd__o21ai_2 _12396_ (.A1(_06593_),
    .A2(_06595_),
    .B1(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__nor2_2 _12397_ (.A(_06628_),
    .B(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__a211o_1 _12398_ (.A1(_06628_),
    .A2(_06630_),
    .B1(_06586_),
    .C1(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__o2111ai_4 _12399_ (.A1(_06608_),
    .A2(_06616_),
    .B1(_06620_),
    .C1(_06624_),
    .D1(_06632_),
    .Y(_00363_));
 sky130_fd_sc_hd__or2_2 _12400_ (.A(_00169_),
    .B(_06584_),
    .X(_00255_));
 sky130_fd_sc_hd__buf_1 _12401_ (.A(_06626_),
    .X(_06633_));
 sky130_fd_sc_hd__inv_2 _12402_ (.A(\e1.alu1.a[27] ),
    .Y(_06634_));
 sky130_fd_sc_hd__buf_1 _12403_ (.A(\e1.alu1.a1.b[27] ),
    .X(_06635_));
 sky130_fd_sc_hd__inv_2 _12404_ (.A(\e1.alu1.a1.b[27] ),
    .Y(_06636_));
 sky130_fd_sc_hd__o22a_2 _12405_ (.A1(_06635_),
    .A2(_06541_),
    .B1(_06636_),
    .B2(_06543_),
    .X(_06637_));
 sky130_fd_sc_hd__buf_1 _12406_ (.A(\e1.alu1.a[27] ),
    .X(_06638_));
 sky130_fd_sc_hd__inv_2 _12407_ (.A(_06637_),
    .Y(_06639_));
 sky130_fd_sc_hd__o22a_2 _12408_ (.A1(_06634_),
    .A2(_06637_),
    .B1(_06638_),
    .B2(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__inv_2 _12409_ (.A(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__nor2_1 _12410_ (.A(_06633_),
    .B(_06631_),
    .Y(_06642_));
 sky130_fd_sc_hd__o32a_1 _12411_ (.A1(_06633_),
    .A2(_06631_),
    .A3(_06641_),
    .B1(_06640_),
    .B2(_06642_),
    .X(_06643_));
 sky130_fd_sc_hd__buf_1 _12412_ (.A(_06638_),
    .X(_06644_));
 sky130_fd_sc_hd__o21ai_2 _12413_ (.A1(_06635_),
    .A2(_06644_),
    .B1(_06598_),
    .Y(_06645_));
 sky130_fd_sc_hd__buf_1 _12414_ (.A(_06636_),
    .X(_06646_));
 sky130_fd_sc_hd__buf_4 _12415_ (.A(_06634_),
    .X(_00081_));
 sky130_fd_sc_hd__buf_1 _12416_ (.A(_06601_),
    .X(_06647_));
 sky130_fd_sc_hd__buf_1 _12417_ (.A(_06580_),
    .X(_06648_));
 sky130_fd_sc_hd__o32a_1 _12418_ (.A1(_06646_),
    .A2(_00081_),
    .A3(_06647_),
    .B1(_00368_),
    .B2(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__o22a_1 _12419_ (.A1(_06635_),
    .A2(_06638_),
    .B1(_06646_),
    .B2(_06634_),
    .X(_06650_));
 sky130_fd_sc_hd__inv_2 _12420_ (.A(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__o22a_1 _12421_ (.A1(_06605_),
    .A2(_00255_),
    .B1(_06608_),
    .B2(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__o2111ai_4 _12422_ (.A1(_06587_),
    .A2(_06643_),
    .B1(_06645_),
    .C1(_06649_),
    .D1(_06652_),
    .Y(_00369_));
 sky130_fd_sc_hd__buf_1 _12423_ (.A(net9),
    .X(_06653_));
 sky130_fd_sc_hd__or2_1 _12424_ (.A(_06653_),
    .B(_00090_),
    .X(_00180_));
 sky130_fd_sc_hd__or2_1 _12425_ (.A(_06564_),
    .B(_00180_),
    .X(_00264_));
 sky130_fd_sc_hd__inv_2 _12426_ (.A(_06552_),
    .Y(_06654_));
 sky130_fd_sc_hd__clkbuf_2 _12427_ (.A(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__buf_2 _12428_ (.A(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__o21ai_2 _12429_ (.A1(_06644_),
    .A2(_06639_),
    .B1(_06633_),
    .Y(_06657_));
 sky130_fd_sc_hd__o2111ai_4 _12430_ (.A1(_06546_),
    .A2(_06593_),
    .B1(_06629_),
    .C1(_06627_),
    .D1(_06640_),
    .Y(_06658_));
 sky130_fd_sc_hd__or2_1 _12431_ (.A(_06547_),
    .B(_06594_),
    .X(_06659_));
 sky130_fd_sc_hd__or4_4 _12432_ (.A(_06628_),
    .B(_06641_),
    .C(_06659_),
    .D(_06539_),
    .X(_06660_));
 sky130_fd_sc_hd__o2111ai_4 _12433_ (.A1(_00081_),
    .A2(_06637_),
    .B1(_06657_),
    .C1(_06658_),
    .D1(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__inv_2 _12434_ (.A(\e1.alu1.a[28] ),
    .Y(_06662_));
 sky130_fd_sc_hd__buf_2 _12435_ (.A(_06662_),
    .X(_00084_));
 sky130_fd_sc_hd__inv_2 _12436_ (.A(\e1.alu1.a1.b[28] ),
    .Y(_06663_));
 sky130_fd_sc_hd__buf_1 _12437_ (.A(_06544_),
    .X(_06664_));
 sky130_fd_sc_hd__o22a_1 _12438_ (.A1(\e1.alu1.a1.b[28] ),
    .A2(_06585_),
    .B1(_06663_),
    .B2(_06664_),
    .X(_06665_));
 sky130_fd_sc_hd__buf_1 _12439_ (.A(\e1.alu1.a[28] ),
    .X(_06666_));
 sky130_fd_sc_hd__inv_2 _12440_ (.A(_06665_),
    .Y(_06667_));
 sky130_fd_sc_hd__o22a_1 _12441_ (.A1(_00084_),
    .A2(_06665_),
    .B1(_06666_),
    .B2(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__or2_1 _12442_ (.A(_06661_),
    .B(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__nand2_1 _12443_ (.A(_06661_),
    .B(_06668_),
    .Y(_06670_));
 sky130_fd_sc_hd__nor2_1 _12444_ (.A(\e1.alu1.a1.b[28] ),
    .B(\e1.alu1.a[28] ),
    .Y(_06671_));
 sky130_fd_sc_hd__clkbuf_2 _12445_ (.A(_06606_),
    .X(_06672_));
 sky130_fd_sc_hd__or2_1 _12446_ (.A(_06663_),
    .B(_06662_),
    .X(_06673_));
 sky130_fd_sc_hd__inv_2 _12447_ (.A(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__clkbuf_2 _12448_ (.A(_06304_),
    .X(_06675_));
 sky130_fd_sc_hd__o21a_1 _12449_ (.A1(_06672_),
    .A2(_06674_),
    .B1(_06675_),
    .X(_06676_));
 sky130_fd_sc_hd__buf_1 _12450_ (.A(_06601_),
    .X(_06677_));
 sky130_fd_sc_hd__buf_1 _12451_ (.A(_06617_),
    .X(_06678_));
 sky130_fd_sc_hd__or2_1 _12452_ (.A(_06561_),
    .B(_00264_),
    .X(_06679_));
 sky130_fd_sc_hd__o221a_1 _12453_ (.A1(_06677_),
    .A2(_06673_),
    .B1(_00374_),
    .B2(_06678_),
    .C1(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__o21ai_1 _12454_ (.A1(_06671_),
    .A2(_06676_),
    .B1(_06680_),
    .Y(_06681_));
 sky130_fd_sc_hd__a31o_1 _12455_ (.A1(_06656_),
    .A2(_06669_),
    .A3(_06670_),
    .B1(_06681_),
    .X(_00375_));
 sky130_fd_sc_hd__buf_1 _12456_ (.A(_06564_),
    .X(_06682_));
 sky130_fd_sc_hd__buf_1 _12457_ (.A(_06653_),
    .X(_06683_));
 sky130_fd_sc_hd__or2_1 _12458_ (.A(_06683_),
    .B(_00127_),
    .X(_00193_));
 sky130_fd_sc_hd__or2_1 _12459_ (.A(_06682_),
    .B(_00193_),
    .X(_00273_));
 sky130_fd_sc_hd__buf_2 _12460_ (.A(_06555_),
    .X(_06684_));
 sky130_fd_sc_hd__inv_2 _12461_ (.A(\e1.alu1.a[29] ),
    .Y(_06685_));
 sky130_fd_sc_hd__clkbuf_2 _12462_ (.A(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__buf_1 _12463_ (.A(\e1.alu1.a1.b[29] ),
    .X(_06687_));
 sky130_fd_sc_hd__inv_2 _12464_ (.A(\e1.alu1.a1.b[29] ),
    .Y(_06688_));
 sky130_fd_sc_hd__o22a_2 _12465_ (.A1(_06687_),
    .A2(_00134_),
    .B1(_06688_),
    .B2(_06664_),
    .X(_06689_));
 sky130_fd_sc_hd__nor2_2 _12466_ (.A(_06685_),
    .B(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__a21oi_4 _12467_ (.A1(_06686_),
    .A2(_06689_),
    .B1(_06690_),
    .Y(_06691_));
 sky130_fd_sc_hd__o21a_1 _12468_ (.A1(_00084_),
    .A2(_06665_),
    .B1(_06670_),
    .X(_06692_));
 sky130_fd_sc_hd__a2bb2oi_2 _12469_ (.A1_N(_06691_),
    .A2_N(_06692_),
    .B1(_06691_),
    .B2(_06692_),
    .Y(_06693_));
 sky130_fd_sc_hd__buf_1 _12470_ (.A(\e1.alu1.a[29] ),
    .X(_06694_));
 sky130_fd_sc_hd__buf_1 _12471_ (.A(_06306_),
    .X(_06695_));
 sky130_fd_sc_hd__clkbuf_2 _12472_ (.A(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__buf_1 _12473_ (.A(_06688_),
    .X(_06697_));
 sky130_fd_sc_hd__clkbuf_4 _12474_ (.A(_06686_),
    .X(_00085_));
 sky130_fd_sc_hd__clkbuf_2 _12475_ (.A(_06569_),
    .X(_06698_));
 sky130_fd_sc_hd__o21a_1 _12476_ (.A1(_06697_),
    .A2(_00085_),
    .B1(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__o22ai_1 _12477_ (.A1(_06687_),
    .A2(_06694_),
    .B1(_06696_),
    .B2(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__buf_1 _12478_ (.A(_06574_),
    .X(_06701_));
 sky130_fd_sc_hd__buf_1 _12479_ (.A(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__or3_2 _12480_ (.A(_06697_),
    .B(_00085_),
    .C(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__o221a_1 _12481_ (.A1(_00380_),
    .A2(_06678_),
    .B1(_06623_),
    .B2(_00273_),
    .C1(_06703_),
    .X(_06704_));
 sky130_fd_sc_hd__o211ai_2 _12482_ (.A1(_06684_),
    .A2(_06693_),
    .B1(_06700_),
    .C1(_06704_),
    .Y(_00381_));
 sky130_fd_sc_hd__clkbuf_1 _12483_ (.A(_06583_),
    .X(_06705_));
 sky130_fd_sc_hd__clkbuf_1 _12484_ (.A(_06683_),
    .X(_06706_));
 sky130_fd_sc_hd__buf_1 _12485_ (.A(\e1.alu1.a1.b[1] ),
    .X(_06707_));
 sky130_fd_sc_hd__clkbuf_2 _12486_ (.A(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__or2_1 _12487_ (.A(_06708_),
    .B(_00089_),
    .X(_00148_));
 sky130_fd_sc_hd__or2_1 _12488_ (.A(_06706_),
    .B(_00148_),
    .X(_00206_));
 sky130_fd_sc_hd__or2_2 _12489_ (.A(_06705_),
    .B(_00206_),
    .X(_00282_));
 sky130_fd_sc_hd__inv_2 _12490_ (.A(\e1.alu1.a[30] ),
    .Y(_06709_));
 sky130_fd_sc_hd__buf_1 _12491_ (.A(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__clkbuf_4 _12492_ (.A(_06710_),
    .X(_00087_));
 sky130_fd_sc_hd__clkbuf_4 _12493_ (.A(_06581_),
    .X(_06711_));
 sky130_fd_sc_hd__inv_2 _12494_ (.A(\e1.alu1.a1.b[30] ),
    .Y(_06712_));
 sky130_fd_sc_hd__buf_1 _12495_ (.A(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__buf_1 _12496_ (.A(_06604_),
    .X(_06714_));
 sky130_fd_sc_hd__o32a_1 _12497_ (.A1(_06713_),
    .A2(_00087_),
    .A3(_06577_),
    .B1(_06714_),
    .B2(_00282_),
    .X(_06715_));
 sky130_fd_sc_hd__clkbuf_2 _12498_ (.A(\e1.alu1.a1.b[30] ),
    .X(_06716_));
 sky130_fd_sc_hd__clkbuf_2 _12499_ (.A(\e1.alu1.a[30] ),
    .X(_06717_));
 sky130_fd_sc_hd__buf_1 _12500_ (.A(_06306_),
    .X(_06718_));
 sky130_fd_sc_hd__buf_2 _12501_ (.A(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__buf_1 _12502_ (.A(_06568_),
    .X(_06720_));
 sky130_fd_sc_hd__o21a_1 _12503_ (.A1(_06713_),
    .A2(_00087_),
    .B1(_06720_),
    .X(_06721_));
 sky130_fd_sc_hd__o22ai_4 _12504_ (.A1(_06716_),
    .A2(_06717_),
    .B1(_06719_),
    .B2(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__buf_1 _12505_ (.A(_06664_),
    .X(_06723_));
 sky130_fd_sc_hd__o22a_1 _12506_ (.A1(_06716_),
    .A2(_00134_),
    .B1(_06712_),
    .B2(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__inv_2 _12507_ (.A(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__o22a_1 _12508_ (.A1(_06710_),
    .A2(_06724_),
    .B1(_06717_),
    .B2(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__nand2_1 _12509_ (.A(_06686_),
    .B(_06689_),
    .Y(_06727_));
 sky130_fd_sc_hd__a31o_1 _12510_ (.A1(_06666_),
    .A2(_06667_),
    .A3(_06727_),
    .B1(_06690_),
    .X(_06728_));
 sky130_fd_sc_hd__a31o_1 _12511_ (.A1(_06668_),
    .A2(_06691_),
    .A3(_06661_),
    .B1(_06728_),
    .X(_06729_));
 sky130_fd_sc_hd__clkbuf_4 _12512_ (.A(_06654_),
    .X(_06730_));
 sky130_fd_sc_hd__nand2_1 _12513_ (.A(_06726_),
    .B(_06729_),
    .Y(_06731_));
 sky130_fd_sc_hd__o211ai_2 _12514_ (.A1(_06726_),
    .A2(_06729_),
    .B1(_06730_),
    .C1(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__o2111ai_4 _12515_ (.A1(_00386_),
    .A2(_06711_),
    .B1(_06715_),
    .C1(_06722_),
    .D1(_06732_),
    .Y(_00387_));
 sky130_fd_sc_hd__inv_2 _12516_ (.A(\e1.alu1.a[31] ),
    .Y(_06733_));
 sky130_fd_sc_hd__buf_1 _12517_ (.A(\e1.alu1.a1.b[0] ),
    .X(_06734_));
 sky130_fd_sc_hd__or2_2 _12518_ (.A(_06733_),
    .B(_06734_),
    .X(_00126_));
 sky130_fd_sc_hd__or2_1 _12519_ (.A(_06707_),
    .B(_00126_),
    .X(_00168_));
 sky130_fd_sc_hd__or2_1 _12520_ (.A(_06706_),
    .B(_00168_),
    .X(_00219_));
 sky130_fd_sc_hd__or2_1 _12521_ (.A(_06705_),
    .B(_00219_),
    .X(_00291_));
 sky130_fd_sc_hd__buf_1 _12522_ (.A(_06733_),
    .X(_00088_));
 sky130_fd_sc_hd__inv_2 _12523_ (.A(\e1.alu1.a1.b[31] ),
    .Y(_06735_));
 sky130_fd_sc_hd__buf_1 _12524_ (.A(_06735_),
    .X(_06736_));
 sky130_fd_sc_hd__o32a_1 _12525_ (.A1(_06736_),
    .A2(_00088_),
    .A3(_06577_),
    .B1(_06714_),
    .B2(_00291_),
    .X(_06737_));
 sky130_fd_sc_hd__clkbuf_2 _12526_ (.A(\e1.alu1.a[31] ),
    .X(_06738_));
 sky130_fd_sc_hd__o21a_1 _12527_ (.A1(_06736_),
    .A2(_00088_),
    .B1(_06720_),
    .X(_06739_));
 sky130_fd_sc_hd__o22ai_4 _12528_ (.A1(\e1.alu1.a1.b[31] ),
    .A2(_06738_),
    .B1(_06719_),
    .B2(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__o21ai_2 _12529_ (.A1(_06710_),
    .A2(_06724_),
    .B1(_06731_),
    .Y(_06741_));
 sky130_fd_sc_hd__inv_2 _12530_ (.A(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__o22a_1 _12531_ (.A1(_06735_),
    .A2(_06733_),
    .B1(\e1.alu1.a1.b[31] ),
    .B2(\e1.alu1.a[31] ),
    .X(_06743_));
 sky130_fd_sc_hd__clkbuf_1 _12532_ (.A(_06743_),
    .X(_06744_));
 sky130_fd_sc_hd__a2bb2o_1 _12533_ (.A1_N(_06723_),
    .A2_N(_06744_),
    .B1(_06723_),
    .B2(_06744_),
    .X(_06745_));
 sky130_fd_sc_hd__inv_2 _12534_ (.A(_06745_),
    .Y(_06746_));
 sky130_fd_sc_hd__clkbuf_2 _12535_ (.A(_06553_),
    .X(_06747_));
 sky130_fd_sc_hd__a221o_1 _12536_ (.A1(_06742_),
    .A2(_06745_),
    .B1(_06741_),
    .B2(_06746_),
    .C1(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__o2111ai_4 _12537_ (.A1(_00392_),
    .A2(_06711_),
    .B1(_06737_),
    .C1(_06740_),
    .D1(_06748_),
    .Y(_00393_));
 sky130_fd_sc_hd__or4_4 _12538_ (.A(\c1.instruction3[3] ),
    .B(\c1.instruction3[2] ),
    .C(\c1.instruction3[4] ),
    .D(\c1.instruction3[6] ),
    .X(_06749_));
 sky130_fd_sc_hd__and3b_1 _12539_ (.A_N(_06749_),
    .B(\c1.instruction3[0] ),
    .C(\c1.instruction3[1] ),
    .X(_06750_));
 sky130_fd_sc_hd__nor2b_4 _12540_ (.A(\c1.instruction3[5] ),
    .B_N(_06750_),
    .Y(ren));
 sky130_fd_sc_hd__and2_2 _12541_ (.A(\c1.instruction3[5] ),
    .B(_06750_),
    .X(wen));
 sky130_fd_sc_hd__inv_2 _12542_ (.A(\c1.instruction3[12] ),
    .Y(_06751_));
 sky130_fd_sc_hd__buf_1 _12543_ (.A(\c1.instruction3[13] ),
    .X(_06752_));
 sky130_fd_sc_hd__inv_2 _12544_ (.A(\c1.instruction3[14] ),
    .Y(_06753_));
 sky130_fd_sc_hd__and3_1 _12545_ (.A(_06751_),
    .B(_06752_),
    .C(_06753_),
    .X(_06754_));
 sky130_fd_sc_hd__buf_1 _12546_ (.A(_06754_),
    .X(_06755_));
 sky130_fd_sc_hd__buf_1 _12547_ (.A(data_address[1]),
    .X(_06756_));
 sky130_fd_sc_hd__o21a_1 _12548_ (.A1(_06751_),
    .A2(_06752_),
    .B1(data_address[0]),
    .X(_06757_));
 sky130_fd_sc_hd__nor2_1 _12549_ (.A(_06756_),
    .B(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__inv_2 _12550_ (.A(\c1.instruction3[13] ),
    .Y(_06759_));
 sky130_fd_sc_hd__nor2_1 _12551_ (.A(_06752_),
    .B(\c1.instruction3[5] ),
    .Y(_06760_));
 sky130_fd_sc_hd__o221a_1 _12552_ (.A1(_06751_),
    .A2(_06759_),
    .B1(_06753_),
    .B2(_06760_),
    .C1(_06750_),
    .X(_06761_));
 sky130_fd_sc_hd__buf_1 _12553_ (.A(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__o21a_2 _12554_ (.A1(_06755_),
    .A2(_06758_),
    .B1(_06762_),
    .X(wstrobe[0]));
 sky130_fd_sc_hd__a21oi_1 _12555_ (.A1(\c1.instruction3[12] ),
    .A2(_06759_),
    .B1(data_address[0]),
    .Y(_06763_));
 sky130_fd_sc_hd__nor2_1 _12556_ (.A(_06756_),
    .B(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__o21a_2 _12557_ (.A1(_06755_),
    .A2(_06764_),
    .B1(_06762_),
    .X(wstrobe[1]));
 sky130_fd_sc_hd__inv_2 _12558_ (.A(data_address[1]),
    .Y(_06765_));
 sky130_fd_sc_hd__nor2_1 _12559_ (.A(_06765_),
    .B(_06757_),
    .Y(_06766_));
 sky130_fd_sc_hd__o21a_4 _12560_ (.A1(_06755_),
    .A2(_06766_),
    .B1(_06762_),
    .X(wstrobe[2]));
 sky130_fd_sc_hd__nor2_1 _12561_ (.A(_06765_),
    .B(_06763_),
    .Y(_06767_));
 sky130_fd_sc_hd__o21a_2 _12562_ (.A1(_06754_),
    .A2(_06767_),
    .B1(_06761_),
    .X(wstrobe[3]));
 sky130_fd_sc_hd__and3_2 _12563_ (.A(_03900_),
    .B(\c1.instruction1[12] ),
    .C(_03897_),
    .X(_00394_));
 sky130_fd_sc_hd__or4_4 _12564_ (.A(\c1.instruction1[28] ),
    .B(\c1.instruction1[27] ),
    .C(\c1.instruction1[26] ),
    .D(\c1.instruction1[25] ),
    .X(_06768_));
 sky130_fd_sc_hd__or3_4 _12565_ (.A(\c1.instruction1[31] ),
    .B(\c1.instruction1[29] ),
    .C(_06768_),
    .X(_06769_));
 sky130_fd_sc_hd__o21a_1 _12566_ (.A1(_03897_),
    .A2(_06769_),
    .B1(_03795_),
    .X(_06770_));
 sky130_fd_sc_hd__buf_1 _12567_ (.A(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__nor2_1 _12568_ (.A(_03858_),
    .B(_06771_),
    .Y(_00395_));
 sky130_fd_sc_hd__buf_1 _12569_ (.A(_03851_),
    .X(_00397_));
 sky130_fd_sc_hd__or2_1 _12570_ (.A(_00397_),
    .B(_06771_),
    .X(_00398_));
 sky130_fd_sc_hd__buf_1 _12571_ (.A(_03846_),
    .X(_00400_));
 sky130_fd_sc_hd__or2_1 _12572_ (.A(_00400_),
    .B(_06771_),
    .X(_00401_));
 sky130_fd_sc_hd__or2_1 _12573_ (.A(_00403_),
    .B(_06770_),
    .X(_00404_));
 sky130_fd_sc_hd__buf_1 _12574_ (.A(_03836_),
    .X(_00406_));
 sky130_fd_sc_hd__or2_1 _12575_ (.A(_00406_),
    .B(_06770_),
    .X(_00407_));
 sky130_fd_sc_hd__a31oi_4 _12576_ (.A1(\c1.instruction1[14] ),
    .A2(_03795_),
    .A3(_06769_),
    .B1(_03792_),
    .Y(_00420_));
 sky130_fd_sc_hd__clkbuf_4 _12577_ (.A(_06309_),
    .X(_00072_));
 sky130_fd_sc_hd__clkbuf_4 _12578_ (.A(_06586_),
    .X(_06772_));
 sky130_fd_sc_hd__buf_1 _12579_ (.A(_06355_),
    .X(_06773_));
 sky130_fd_sc_hd__buf_1 _12580_ (.A(_06343_),
    .X(_06774_));
 sky130_fd_sc_hd__buf_1 _12581_ (.A(_06526_),
    .X(_06775_));
 sky130_fd_sc_hd__o21ai_1 _12582_ (.A1(_06775_),
    .A2(_06388_),
    .B1(_06535_),
    .Y(_06776_));
 sky130_fd_sc_hd__a31o_1 _12583_ (.A1(_06773_),
    .A2(_06774_),
    .A3(_06776_),
    .B1(_06528_),
    .X(_06777_));
 sky130_fd_sc_hd__and2_1 _12584_ (.A(_06322_),
    .B(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__inv_2 _12585_ (.A(_06333_),
    .Y(_06779_));
 sky130_fd_sc_hd__nor2_1 _12586_ (.A(_06321_),
    .B(_06778_),
    .Y(_06780_));
 sky130_fd_sc_hd__o32a_2 _12587_ (.A1(_06321_),
    .A2(_06778_),
    .A3(_06779_),
    .B1(_06333_),
    .B2(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__buf_1 _12588_ (.A(_06323_),
    .X(_06782_));
 sky130_fd_sc_hd__o21ai_2 _12589_ (.A1(_06782_),
    .A2(_06324_),
    .B1(_06598_),
    .Y(_06783_));
 sky130_fd_sc_hd__buf_4 _12590_ (.A(_06536_),
    .X(_00073_));
 sky130_fd_sc_hd__buf_1 _12591_ (.A(_06328_),
    .X(_06784_));
 sky130_fd_sc_hd__o32a_1 _12592_ (.A1(_00073_),
    .A2(_06784_),
    .A3(_06647_),
    .B1(_00344_),
    .B2(_06648_),
    .X(_06785_));
 sky130_fd_sc_hd__buf_1 _12593_ (.A(_06672_),
    .X(_06786_));
 sky130_fd_sc_hd__o22a_1 _12594_ (.A1(_06782_),
    .A2(_06324_),
    .B1(_00073_),
    .B2(_06784_),
    .X(_06787_));
 sky130_fd_sc_hd__inv_2 _12595_ (.A(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__o22a_1 _12596_ (.A1(_00220_),
    .A2(_06605_),
    .B1(_06786_),
    .B2(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__o2111ai_4 _12597_ (.A1(_06772_),
    .A2(_06781_),
    .B1(_06783_),
    .C1(_06785_),
    .D1(_06789_),
    .Y(_00345_));
 sky130_fd_sc_hd__nor2_1 _12598_ (.A(_06322_),
    .B(_06777_),
    .Y(_06790_));
 sky130_fd_sc_hd__buf_1 _12599_ (.A(_06315_),
    .X(_06791_));
 sky130_fd_sc_hd__buf_1 _12600_ (.A(_06575_),
    .X(_06792_));
 sky130_fd_sc_hd__o32a_1 _12601_ (.A1(_06791_),
    .A2(_00072_),
    .A3(_06792_),
    .B1(_00207_),
    .B2(_06562_),
    .X(_06793_));
 sky130_fd_sc_hd__buf_1 _12602_ (.A(\e1.alu1.a[22] ),
    .X(_06794_));
 sky130_fd_sc_hd__o22a_1 _12603_ (.A1(_06791_),
    .A2(_00072_),
    .B1(_06310_),
    .B2(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__inv_2 _12604_ (.A(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__buf_1 _12605_ (.A(_06305_),
    .X(_06797_));
 sky130_fd_sc_hd__o21ai_1 _12606_ (.A1(_06310_),
    .A2(_06794_),
    .B1(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__o221a_1 _12607_ (.A1(_06607_),
    .A2(_06796_),
    .B1(_00338_),
    .B2(_06580_),
    .C1(_06798_),
    .X(_06799_));
 sky130_fd_sc_hd__o311a_1 _12608_ (.A1(_06747_),
    .A2(_06778_),
    .A3(_06790_),
    .B1(_06793_),
    .C1(_06799_),
    .X(_06800_));
 sky130_fd_sc_hd__inv_2 _12609_ (.A(_06800_),
    .Y(_00339_));
 sky130_fd_sc_hd__buf_4 _12610_ (.A(_06345_),
    .X(_00070_));
 sky130_fd_sc_hd__clkbuf_4 _12611_ (.A(_06335_),
    .X(_00069_));
 sky130_fd_sc_hd__nand2_1 _12612_ (.A(_06774_),
    .B(_06776_),
    .Y(_06801_));
 sky130_fd_sc_hd__o21a_1 _12613_ (.A1(_00069_),
    .A2(_06340_),
    .B1(_06801_),
    .X(_06802_));
 sky130_fd_sc_hd__a2bb2oi_2 _12614_ (.A1_N(_06773_),
    .A2_N(_06802_),
    .B1(_06773_),
    .B2(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__buf_1 _12615_ (.A(\e1.alu1.a[21] ),
    .X(_06804_));
 sky130_fd_sc_hd__clkbuf_2 _12616_ (.A(_06695_),
    .X(_06805_));
 sky130_fd_sc_hd__o21ai_2 _12617_ (.A1(_06804_),
    .A2(_06346_),
    .B1(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__buf_1 _12618_ (.A(_06349_),
    .X(_06807_));
 sky130_fd_sc_hd__o32a_2 _12619_ (.A1(_00070_),
    .A2(_06807_),
    .A3(_06647_),
    .B1(_00332_),
    .B2(_06648_),
    .X(_06808_));
 sky130_fd_sc_hd__buf_1 _12620_ (.A(_06604_),
    .X(_06809_));
 sky130_fd_sc_hd__o22a_1 _12621_ (.A1(_06804_),
    .A2(_06346_),
    .B1(_00070_),
    .B2(_06807_),
    .X(_06810_));
 sky130_fd_sc_hd__inv_2 _12622_ (.A(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__o22a_1 _12623_ (.A1(_00194_),
    .A2(_06809_),
    .B1(_06786_),
    .B2(_06811_),
    .X(_06812_));
 sky130_fd_sc_hd__o2111ai_4 _12624_ (.A1(_06772_),
    .A2(_06803_),
    .B1(_06806_),
    .C1(_06808_),
    .D1(_06812_),
    .Y(_00333_));
 sky130_fd_sc_hd__or2_1 _12625_ (.A(_06774_),
    .B(_06776_),
    .X(_06813_));
 sky130_fd_sc_hd__buf_1 _12626_ (.A(_06341_),
    .X(_06814_));
 sky130_fd_sc_hd__buf_1 _12627_ (.A(_06338_),
    .X(_06815_));
 sky130_fd_sc_hd__o22a_1 _12628_ (.A1(_06814_),
    .A2(_06336_),
    .B1(_06335_),
    .B2(_06815_),
    .X(_06816_));
 sky130_fd_sc_hd__a2bb2o_1 _12629_ (.A1_N(_00181_),
    .A2_N(_06623_),
    .B1(_06698_),
    .B2(_06816_),
    .X(_06817_));
 sky130_fd_sc_hd__o21ai_1 _12630_ (.A1(_06814_),
    .A2(_06336_),
    .B1(_06307_),
    .Y(_06818_));
 sky130_fd_sc_hd__o32a_1 _12631_ (.A1(_00069_),
    .A2(_06815_),
    .A3(_06792_),
    .B1(_00326_),
    .B2(_06678_),
    .X(_06819_));
 sky130_fd_sc_hd__nand2_1 _12632_ (.A(_06818_),
    .B(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__a311o_1 _12633_ (.A1(_06656_),
    .A2(_06801_),
    .A3(_06813_),
    .B1(_06817_),
    .C1(_06820_),
    .X(_00327_));
 sky130_fd_sc_hd__clkbuf_4 _12634_ (.A(_06357_),
    .X(_00066_));
 sky130_fd_sc_hd__clkbuf_4 _12635_ (.A(_06364_),
    .X(_00065_));
 sky130_fd_sc_hd__buf_1 _12636_ (.A(_06387_),
    .X(_06821_));
 sky130_fd_sc_hd__inv_2 _12637_ (.A(_06526_),
    .Y(_06822_));
 sky130_fd_sc_hd__a31o_1 _12638_ (.A1(_06821_),
    .A2(_06379_),
    .A3(_06822_),
    .B1(_06531_),
    .X(_06823_));
 sky130_fd_sc_hd__and2_1 _12639_ (.A(_06369_),
    .B(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__inv_2 _12640_ (.A(_06363_),
    .Y(_06825_));
 sky130_fd_sc_hd__nor2_1 _12641_ (.A(_06533_),
    .B(_06824_),
    .Y(_06826_));
 sky130_fd_sc_hd__o32a_2 _12642_ (.A1(_06533_),
    .A2(_06824_),
    .A3(_06825_),
    .B1(_06363_),
    .B2(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__buf_1 _12643_ (.A(_06361_),
    .X(_06828_));
 sky130_fd_sc_hd__o21ai_2 _12644_ (.A1(_06828_),
    .A2(_06358_),
    .B1(_06805_),
    .Y(_06829_));
 sky130_fd_sc_hd__buf_1 _12645_ (.A(_06359_),
    .X(_06830_));
 sky130_fd_sc_hd__o32a_1 _12646_ (.A1(_00066_),
    .A2(_06830_),
    .A3(_06677_),
    .B1(_00320_),
    .B2(_06618_),
    .X(_06831_));
 sky130_fd_sc_hd__o22a_1 _12647_ (.A1(_06828_),
    .A2(_06358_),
    .B1(_00066_),
    .B2(_06830_),
    .X(_06832_));
 sky130_fd_sc_hd__inv_2 _12648_ (.A(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__o22a_1 _12649_ (.A1(_00170_),
    .A2(_06809_),
    .B1(_06786_),
    .B2(_06833_),
    .X(_06834_));
 sky130_fd_sc_hd__o2111ai_4 _12650_ (.A1(_06772_),
    .A2(_06827_),
    .B1(_06829_),
    .C1(_06831_),
    .D1(_06834_),
    .Y(_00321_));
 sky130_fd_sc_hd__nor2_1 _12651_ (.A(_06369_),
    .B(_06823_),
    .Y(_06835_));
 sky130_fd_sc_hd__buf_1 _12652_ (.A(_06366_),
    .X(_06836_));
 sky130_fd_sc_hd__o32a_1 _12653_ (.A1(_06836_),
    .A2(_00065_),
    .A3(_06576_),
    .B1(_00150_),
    .B2(_06562_),
    .X(_06837_));
 sky130_fd_sc_hd__buf_1 _12654_ (.A(\e1.alu1.a[18] ),
    .X(_06838_));
 sky130_fd_sc_hd__o22a_1 _12655_ (.A1(_06836_),
    .A2(_00065_),
    .B1(_06365_),
    .B2(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__inv_2 _12656_ (.A(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__o21ai_1 _12657_ (.A1(_06365_),
    .A2(_06838_),
    .B1(_06797_),
    .Y(_06841_));
 sky130_fd_sc_hd__o221a_1 _12658_ (.A1(_06607_),
    .A2(_06840_),
    .B1(_00314_),
    .B2(_06617_),
    .C1(_06841_),
    .X(_06842_));
 sky130_fd_sc_hd__o311a_1 _12659_ (.A1(_06747_),
    .A2(_06824_),
    .A3(_06835_),
    .B1(_06837_),
    .C1(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__inv_2 _12660_ (.A(_06843_),
    .Y(_00315_));
 sky130_fd_sc_hd__buf_1 _12661_ (.A(_06371_),
    .X(_06844_));
 sky130_fd_sc_hd__clkbuf_4 _12662_ (.A(_06844_),
    .X(_00062_));
 sky130_fd_sc_hd__buf_2 _12663_ (.A(_06554_),
    .X(_06845_));
 sky130_fd_sc_hd__o22a_1 _12664_ (.A1(_06844_),
    .A2(_06376_),
    .B1(_06775_),
    .B2(_06380_),
    .X(_06846_));
 sky130_fd_sc_hd__a2bb2oi_2 _12665_ (.A1_N(_06821_),
    .A2_N(_06846_),
    .B1(_06821_),
    .B2(_06846_),
    .Y(_06847_));
 sky130_fd_sc_hd__buf_1 _12666_ (.A(\e1.alu1.a[17] ),
    .X(_06848_));
 sky130_fd_sc_hd__o21ai_2 _12667_ (.A1(_06848_),
    .A2(_06383_),
    .B1(_06805_),
    .Y(_06849_));
 sky130_fd_sc_hd__buf_1 _12668_ (.A(_06384_),
    .X(_06850_));
 sky130_fd_sc_hd__o32a_1 _12669_ (.A1(_00063_),
    .A2(_06850_),
    .A3(_06677_),
    .B1(_00308_),
    .B2(_06618_),
    .X(_06851_));
 sky130_fd_sc_hd__buf_1 _12670_ (.A(_06606_),
    .X(_06852_));
 sky130_fd_sc_hd__o22a_1 _12671_ (.A1(_06848_),
    .A2(_06383_),
    .B1(_06382_),
    .B2(_06850_),
    .X(_06853_));
 sky130_fd_sc_hd__inv_2 _12672_ (.A(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__o22a_1 _12673_ (.A1(_00129_),
    .A2(_06809_),
    .B1(_06852_),
    .B2(_06854_),
    .X(_06855_));
 sky130_fd_sc_hd__o2111ai_4 _12674_ (.A1(_06845_),
    .A2(_06847_),
    .B1(_06849_),
    .C1(_06851_),
    .D1(_06855_),
    .Y(_00309_));
 sky130_fd_sc_hd__buf_1 _12675_ (.A(_06372_),
    .X(_06856_));
 sky130_fd_sc_hd__buf_1 _12676_ (.A(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__buf_1 _12677_ (.A(_06702_),
    .X(_06858_));
 sky130_fd_sc_hd__o32a_1 _12678_ (.A1(_00062_),
    .A2(_06857_),
    .A3(_06858_),
    .B1(_00092_),
    .B2(_06714_),
    .X(_06859_));
 sky130_fd_sc_hd__o21ai_1 _12679_ (.A1(_06844_),
    .A2(_06857_),
    .B1(_06720_),
    .Y(_06860_));
 sky130_fd_sc_hd__a22o_1 _12680_ (.A1(_00062_),
    .A2(_06857_),
    .B1(_06619_),
    .B2(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__clkbuf_2 _12681_ (.A(_06553_),
    .X(_06862_));
 sky130_fd_sc_hd__a221o_1 _12682_ (.A1(_06822_),
    .A2(_06379_),
    .B1(_06775_),
    .B2(_06380_),
    .C1(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__o2111ai_4 _12683_ (.A1(_00302_),
    .A2(_06711_),
    .B1(_06859_),
    .C1(_06861_),
    .D1(_06863_),
    .Y(_00303_));
 sky130_fd_sc_hd__buf_1 _12684_ (.A(_06420_),
    .X(_06864_));
 sky130_fd_sc_hd__clkbuf_1 _12685_ (.A(_06413_),
    .X(_06865_));
 sky130_fd_sc_hd__buf_1 _12686_ (.A(_06513_),
    .X(_06866_));
 sky130_fd_sc_hd__o21ai_1 _12687_ (.A1(_06866_),
    .A2(_06453_),
    .B1(_06522_),
    .Y(_06867_));
 sky130_fd_sc_hd__a31o_1 _12688_ (.A1(_06864_),
    .A2(_06865_),
    .A3(_06867_),
    .B1(_06515_),
    .X(_06868_));
 sky130_fd_sc_hd__nand2_2 _12689_ (.A(_06405_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__and2_1 _12690_ (.A(_06404_),
    .B(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__a2bb2oi_2 _12691_ (.A1_N(_06396_),
    .A2_N(_06870_),
    .B1(_06396_),
    .B2(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__buf_1 _12692_ (.A(_06389_),
    .X(_06872_));
 sky130_fd_sc_hd__buf_2 _12693_ (.A(_06523_),
    .X(_00057_));
 sky130_fd_sc_hd__buf_1 _12694_ (.A(_06391_),
    .X(_06873_));
 sky130_fd_sc_hd__o21a_1 _12695_ (.A1(_00057_),
    .A2(_06873_),
    .B1(_06698_),
    .X(_06874_));
 sky130_fd_sc_hd__o22ai_1 _12696_ (.A1(_06872_),
    .A2(_06390_),
    .B1(_06696_),
    .B2(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__buf_1 _12697_ (.A(_06559_),
    .X(_06876_));
 sky130_fd_sc_hd__buf_1 _12698_ (.A(_06876_),
    .X(_06877_));
 sky130_fd_sc_hd__or2_1 _12699_ (.A(_06558_),
    .B(_06579_),
    .X(_06878_));
 sky130_fd_sc_hd__buf_1 _12700_ (.A(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__buf_1 _12701_ (.A(_06879_),
    .X(_06880_));
 sky130_fd_sc_hd__clkbuf_1 _12702_ (.A(_06701_),
    .X(_06881_));
 sky130_fd_sc_hd__or3_2 _12703_ (.A(_00057_),
    .B(_06873_),
    .C(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__o221a_1 _12704_ (.A1(_00292_),
    .A2(_06877_),
    .B1(_00296_),
    .B2(_06880_),
    .C1(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__o211ai_2 _12705_ (.A1(_06684_),
    .A2(_06871_),
    .B1(_06875_),
    .C1(_06883_),
    .Y(_00297_));
 sky130_fd_sc_hd__clkbuf_2 _12706_ (.A(_06879_),
    .X(_06884_));
 sky130_fd_sc_hd__buf_2 _12707_ (.A(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__buf_1 _12708_ (.A(_06402_),
    .X(_06886_));
 sky130_fd_sc_hd__buf_2 _12709_ (.A(_06398_),
    .X(_00056_));
 sky130_fd_sc_hd__buf_1 _12710_ (.A(_06876_),
    .X(_06887_));
 sky130_fd_sc_hd__o32a_1 _12711_ (.A1(_06886_),
    .A2(_00056_),
    .A3(_06858_),
    .B1(_00283_),
    .B2(_06887_),
    .X(_06888_));
 sky130_fd_sc_hd__clkbuf_2 _12712_ (.A(\e1.alu1.a[14] ),
    .X(_06889_));
 sky130_fd_sc_hd__buf_2 _12713_ (.A(_06718_),
    .X(_06890_));
 sky130_fd_sc_hd__buf_1 _12714_ (.A(_06568_),
    .X(_06891_));
 sky130_fd_sc_hd__buf_1 _12715_ (.A(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__o21a_1 _12716_ (.A1(_06886_),
    .A2(_00056_),
    .B1(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__o22ai_4 _12717_ (.A1(_06399_),
    .A2(_06889_),
    .B1(_06890_),
    .B2(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__o211ai_4 _12718_ (.A1(_06405_),
    .A2(_06868_),
    .B1(_06730_),
    .C1(_06869_),
    .Y(_06895_));
 sky130_fd_sc_hd__o2111ai_4 _12719_ (.A1(_00288_),
    .A2(_06885_),
    .B1(_06888_),
    .C1(_06894_),
    .D1(_06895_),
    .Y(_00289_));
 sky130_fd_sc_hd__clkbuf_4 _12720_ (.A(_06407_),
    .X(_00053_));
 sky130_fd_sc_hd__nand2_1 _12721_ (.A(_06865_),
    .B(_06867_),
    .Y(_06896_));
 sky130_fd_sc_hd__o21a_1 _12722_ (.A1(_00053_),
    .A2(_06410_),
    .B1(_06896_),
    .X(_06897_));
 sky130_fd_sc_hd__a2bb2oi_2 _12723_ (.A1_N(_06864_),
    .A2_N(_06897_),
    .B1(_06864_),
    .B2(_06897_),
    .Y(_06898_));
 sky130_fd_sc_hd__buf_1 _12724_ (.A(\e1.alu1.a[13] ),
    .X(_06899_));
 sky130_fd_sc_hd__buf_2 _12725_ (.A(_06415_),
    .X(_00054_));
 sky130_fd_sc_hd__buf_1 _12726_ (.A(_06417_),
    .X(_06900_));
 sky130_fd_sc_hd__buf_1 _12727_ (.A(_06569_),
    .X(_06901_));
 sky130_fd_sc_hd__o21a_1 _12728_ (.A1(_00054_),
    .A2(_06900_),
    .B1(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__o22ai_1 _12729_ (.A1(_06899_),
    .A2(_06416_),
    .B1(_06696_),
    .B2(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__or3_1 _12730_ (.A(_00054_),
    .B(_06900_),
    .C(_06881_),
    .X(_06904_));
 sky130_fd_sc_hd__o221a_1 _12731_ (.A1(_00274_),
    .A2(_06877_),
    .B1(_00279_),
    .B2(_06880_),
    .C1(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__o211ai_2 _12732_ (.A1(_06684_),
    .A2(_06898_),
    .B1(_06903_),
    .C1(_06905_),
    .Y(_00280_));
 sky130_fd_sc_hd__inv_2 _12733_ (.A(_00212_),
    .Y(_00284_));
 sky130_fd_sc_hd__inv_2 _12734_ (.A(_00199_),
    .Y(_00275_));
 sky130_fd_sc_hd__or2_1 _12735_ (.A(_06865_),
    .B(_06867_),
    .X(_06906_));
 sky130_fd_sc_hd__nor2_2 _12736_ (.A(_06411_),
    .B(\e1.alu1.a1.b[12] ),
    .Y(_06907_));
 sky130_fd_sc_hd__nor2_2 _12737_ (.A(_00053_),
    .B(_06409_),
    .Y(_06908_));
 sky130_fd_sc_hd__o21a_1 _12738_ (.A1(_06672_),
    .A2(_06908_),
    .B1(_06675_),
    .X(_06909_));
 sky130_fd_sc_hd__inv_2 _12739_ (.A(_06575_),
    .Y(_06910_));
 sky130_fd_sc_hd__buf_1 _12740_ (.A(_06559_),
    .X(_06911_));
 sky130_fd_sc_hd__buf_1 _12741_ (.A(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__o2bb2a_1 _12742_ (.A1_N(_06910_),
    .A2_N(_06908_),
    .B1(_00265_),
    .B2(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__o221ai_2 _12743_ (.A1(_00270_),
    .A2(_06884_),
    .B1(_06907_),
    .B2(_06909_),
    .C1(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__a31o_1 _12744_ (.A1(_06656_),
    .A2(_06896_),
    .A3(_06906_),
    .B1(_06914_),
    .X(_00271_));
 sky130_fd_sc_hd__buf_1 _12745_ (.A(_06555_),
    .X(_06915_));
 sky130_fd_sc_hd__buf_1 _12746_ (.A(_06452_),
    .X(_06916_));
 sky130_fd_sc_hd__inv_2 _12747_ (.A(_06513_),
    .Y(_06917_));
 sky130_fd_sc_hd__a31o_1 _12748_ (.A1(_06916_),
    .A2(_06444_),
    .A3(_06917_),
    .B1(_06519_),
    .X(_06918_));
 sky130_fd_sc_hd__nand2_2 _12749_ (.A(_06436_),
    .B(_06918_),
    .Y(_06919_));
 sky130_fd_sc_hd__and2_1 _12750_ (.A(_06434_),
    .B(_06919_),
    .X(_06920_));
 sky130_fd_sc_hd__a2bb2oi_1 _12751_ (.A1_N(_06428_),
    .A2_N(_06920_),
    .B1(_06428_),
    .B2(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__buf_1 _12752_ (.A(_06426_),
    .X(_06922_));
 sky130_fd_sc_hd__buf_1 _12753_ (.A(_06718_),
    .X(_06923_));
 sky130_fd_sc_hd__clkbuf_4 _12754_ (.A(_06517_),
    .X(_00050_));
 sky130_fd_sc_hd__buf_1 _12755_ (.A(_06424_),
    .X(_06924_));
 sky130_fd_sc_hd__o21a_1 _12756_ (.A1(_00050_),
    .A2(_06924_),
    .B1(_06901_),
    .X(_06925_));
 sky130_fd_sc_hd__o22ai_1 _12757_ (.A1(_06922_),
    .A2(_06423_),
    .B1(_06923_),
    .B2(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__or3_2 _12758_ (.A(_00050_),
    .B(_06924_),
    .C(_06881_),
    .X(_06927_));
 sky130_fd_sc_hd__o221a_1 _12759_ (.A1(_00256_),
    .A2(_06877_),
    .B1(_00261_),
    .B2(_06880_),
    .C1(_06927_),
    .X(_06928_));
 sky130_fd_sc_hd__o211ai_1 _12760_ (.A1(_06915_),
    .A2(_06921_),
    .B1(_06926_),
    .C1(_06928_),
    .Y(_00262_));
 sky130_fd_sc_hd__inv_2 _12761_ (.A(_00186_),
    .Y(_00266_));
 sky130_fd_sc_hd__clkbuf_4 _12762_ (.A(_06430_),
    .X(_00049_));
 sky130_fd_sc_hd__buf_1 _12763_ (.A(_06432_),
    .X(_06929_));
 sky130_fd_sc_hd__o32a_1 _12764_ (.A1(_00049_),
    .A2(_06929_),
    .A3(_06858_),
    .B1(_00247_),
    .B2(_06887_),
    .X(_06930_));
 sky130_fd_sc_hd__clkbuf_2 _12765_ (.A(\e1.alu1.a[10] ),
    .X(_06931_));
 sky130_fd_sc_hd__o21a_1 _12766_ (.A1(_00049_),
    .A2(_06929_),
    .B1(_06892_),
    .X(_06932_));
 sky130_fd_sc_hd__o22ai_4 _12767_ (.A1(_06931_),
    .A2(_06431_),
    .B1(_06890_),
    .B2(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__o211ai_4 _12768_ (.A1(_06436_),
    .A2(_06918_),
    .B1(_06730_),
    .C1(_06919_),
    .Y(_06934_));
 sky130_fd_sc_hd__o2111ai_4 _12769_ (.A1(_00252_),
    .A2(_06885_),
    .B1(_06930_),
    .C1(_06933_),
    .D1(_06934_),
    .Y(_00253_));
 sky130_fd_sc_hd__or2_1 _12770_ (.A(_06706_),
    .B(_00173_),
    .X(_00257_));
 sky130_fd_sc_hd__buf_1 _12771_ (.A(_06461_),
    .X(_06935_));
 sky130_fd_sc_hd__nand2_1 _12772_ (.A(_06935_),
    .B(_00154_),
    .Y(_00248_));
 sky130_fd_sc_hd__clkbuf_4 _12773_ (.A(_06447_),
    .X(_00047_));
 sky130_fd_sc_hd__buf_1 _12774_ (.A(_06438_),
    .X(_06936_));
 sky130_fd_sc_hd__clkbuf_4 _12775_ (.A(_06936_),
    .X(_00046_));
 sky130_fd_sc_hd__o22a_1 _12776_ (.A1(_06936_),
    .A2(_06441_),
    .B1(_06866_),
    .B2(_06445_),
    .X(_06937_));
 sky130_fd_sc_hd__a2bb2oi_1 _12777_ (.A1_N(_06916_),
    .A2_N(_06937_),
    .B1(_06916_),
    .B2(_06937_),
    .Y(_06938_));
 sky130_fd_sc_hd__buf_1 _12778_ (.A(\e1.alu1.a[9] ),
    .X(_06939_));
 sky130_fd_sc_hd__buf_1 _12779_ (.A(_06449_),
    .X(_06940_));
 sky130_fd_sc_hd__o21a_1 _12780_ (.A1(_00047_),
    .A2(_06940_),
    .B1(_06901_),
    .X(_06941_));
 sky130_fd_sc_hd__o22ai_1 _12781_ (.A1(_06939_),
    .A2(_06448_),
    .B1(_06923_),
    .B2(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__buf_1 _12782_ (.A(_06911_),
    .X(_06943_));
 sky130_fd_sc_hd__buf_1 _12783_ (.A(_06878_),
    .X(_06944_));
 sky130_fd_sc_hd__clkbuf_1 _12784_ (.A(_06701_),
    .X(_06945_));
 sky130_fd_sc_hd__or3_1 _12785_ (.A(_00047_),
    .B(_06940_),
    .C(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__o221a_1 _12786_ (.A1(_00238_),
    .A2(_06943_),
    .B1(_00243_),
    .B2(_06944_),
    .C1(_06946_),
    .X(_06947_));
 sky130_fd_sc_hd__o211ai_1 _12787_ (.A1(_06915_),
    .A2(_06938_),
    .B1(_06942_),
    .C1(_06947_),
    .Y(_00244_));
 sky130_fd_sc_hd__buf_1 _12788_ (.A(_06440_),
    .X(_06948_));
 sky130_fd_sc_hd__buf_1 _12789_ (.A(_06702_),
    .X(_06949_));
 sky130_fd_sc_hd__o32a_1 _12790_ (.A1(_00046_),
    .A2(_06948_),
    .A3(_06949_),
    .B1(_00229_),
    .B2(_06887_),
    .X(_06950_));
 sky130_fd_sc_hd__clkbuf_2 _12791_ (.A(_06442_),
    .X(_06951_));
 sky130_fd_sc_hd__o21a_1 _12792_ (.A1(_00046_),
    .A2(_06948_),
    .B1(_06892_),
    .X(_06952_));
 sky130_fd_sc_hd__o22ai_4 _12793_ (.A1(_06951_),
    .A2(_06439_),
    .B1(_06890_),
    .B2(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__a221o_1 _12794_ (.A1(_06917_),
    .A2(_06444_),
    .B1(_06866_),
    .B2(_06445_),
    .C1(_06862_),
    .X(_06954_));
 sky130_fd_sc_hd__o2111ai_4 _12795_ (.A1(_00234_),
    .A2(_06885_),
    .B1(_06950_),
    .C1(_06953_),
    .D1(_06954_),
    .Y(_00235_));
 sky130_fd_sc_hd__nor2_1 _12796_ (.A(_06708_),
    .B(_00131_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2_1 _12797_ (.A(_06935_),
    .B(_00132_),
    .Y(_00239_));
 sky130_fd_sc_hd__buf_1 _12798_ (.A(_06498_),
    .X(_06955_));
 sky130_fd_sc_hd__clkbuf_2 _12799_ (.A(_06505_),
    .X(_06956_));
 sky130_fd_sc_hd__clkbuf_2 _12800_ (.A(_06475_),
    .X(_06957_));
 sky130_fd_sc_hd__a31o_1 _12801_ (.A1(_06955_),
    .A2(_06956_),
    .A3(_06957_),
    .B1(_06510_),
    .X(_06958_));
 sky130_fd_sc_hd__nand2_2 _12802_ (.A(_06508_),
    .B(_06958_),
    .Y(_06959_));
 sky130_fd_sc_hd__and2_1 _12803_ (.A(_06489_),
    .B(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__a2bb2oi_1 _12804_ (.A1_N(_06507_),
    .A2_N(_06960_),
    .B1(_06507_),
    .B2(_06960_),
    .Y(_06961_));
 sky130_fd_sc_hd__buf_1 _12805_ (.A(_06476_),
    .X(_06962_));
 sky130_fd_sc_hd__buf_4 _12806_ (.A(_06477_),
    .X(_00042_));
 sky130_fd_sc_hd__buf_1 _12807_ (.A(_06479_),
    .X(_06963_));
 sky130_fd_sc_hd__o21a_1 _12808_ (.A1(_00042_),
    .A2(_06963_),
    .B1(_06570_),
    .X(_06964_));
 sky130_fd_sc_hd__o22ai_1 _12809_ (.A1(_06962_),
    .A2(_06478_),
    .B1(_06923_),
    .B2(_06964_),
    .Y(_06965_));
 sky130_fd_sc_hd__buf_1 _12810_ (.A(_06944_),
    .X(_06966_));
 sky130_fd_sc_hd__or2_1 _12811_ (.A(_06682_),
    .B(_00224_),
    .X(_00225_));
 sky130_fd_sc_hd__or3_1 _12812_ (.A(_00042_),
    .B(_06963_),
    .C(_06945_),
    .X(_06967_));
 sky130_fd_sc_hd__o221a_1 _12813_ (.A1(_00221_),
    .A2(_06943_),
    .B1(_06966_),
    .B2(_00225_),
    .C1(_06967_),
    .X(_06968_));
 sky130_fd_sc_hd__o211ai_1 _12814_ (.A1(_06915_),
    .A2(_06961_),
    .B1(_06965_),
    .C1(_06968_),
    .Y(_00226_));
 sky130_fd_sc_hd__buf_1 _12815_ (.A(_06467_),
    .X(_06969_));
 sky130_fd_sc_hd__clkinv_4 _12816_ (.A(\e1.alu1.a[0] ),
    .Y(_00031_));
 sky130_fd_sc_hd__nor2_2 _12817_ (.A(net11),
    .B(_00031_),
    .Y(_00024_));
 sky130_fd_sc_hd__nand2_1 _12818_ (.A(_06969_),
    .B(_00024_),
    .Y(_06970_));
 sky130_fd_sc_hd__or2_1 _12819_ (.A(_06683_),
    .B(_06970_),
    .X(_00230_));
 sky130_fd_sc_hd__buf_4 _12820_ (.A(_06485_),
    .X(_00041_));
 sky130_fd_sc_hd__clkbuf_4 _12821_ (.A(_06966_),
    .X(_06971_));
 sky130_fd_sc_hd__buf_1 _12822_ (.A(_06565_),
    .X(_06972_));
 sky130_fd_sc_hd__or2_1 _12823_ (.A(_00284_),
    .B(_06972_),
    .X(_06973_));
 sky130_fd_sc_hd__clkbuf_2 _12824_ (.A(_06973_),
    .X(_00213_));
 sky130_fd_sc_hd__buf_1 _12825_ (.A(_06487_),
    .X(_06974_));
 sky130_fd_sc_hd__buf_1 _12826_ (.A(_06876_),
    .X(_06975_));
 sky130_fd_sc_hd__o32a_1 _12827_ (.A1(_00041_),
    .A2(_06974_),
    .A3(_06949_),
    .B1(_00208_),
    .B2(_06975_),
    .X(_06976_));
 sky130_fd_sc_hd__clkbuf_2 _12828_ (.A(\e1.alu1.a[6] ),
    .X(_06977_));
 sky130_fd_sc_hd__clkbuf_4 _12829_ (.A(_06797_),
    .X(_06978_));
 sky130_fd_sc_hd__buf_1 _12830_ (.A(_06891_),
    .X(_06979_));
 sky130_fd_sc_hd__o21a_1 _12831_ (.A1(_00041_),
    .A2(_06974_),
    .B1(_06979_),
    .X(_06980_));
 sky130_fd_sc_hd__o22ai_4 _12832_ (.A1(_06977_),
    .A2(_06486_),
    .B1(_06978_),
    .B2(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__o211ai_4 _12833_ (.A1(_06508_),
    .A2(_06958_),
    .B1(_06655_),
    .C1(_06959_),
    .Y(_06982_));
 sky130_fd_sc_hd__o2111ai_4 _12834_ (.A1(_06971_),
    .A2(_00213_),
    .B1(_06976_),
    .C1(_06981_),
    .D1(_06982_),
    .Y(_00214_));
 sky130_fd_sc_hd__inv_2 _12835_ (.A(_00210_),
    .Y(_00211_));
 sky130_fd_sc_hd__buf_4 _12836_ (.A(_06493_),
    .X(_00039_));
 sky130_fd_sc_hd__buf_1 _12837_ (.A(_06499_),
    .X(_06983_));
 sky130_fd_sc_hd__clkbuf_4 _12838_ (.A(_06983_),
    .X(_00038_));
 sky130_fd_sc_hd__nand2_2 _12839_ (.A(_06957_),
    .B(_06956_),
    .Y(_06984_));
 sky130_fd_sc_hd__o21a_1 _12840_ (.A1(_06983_),
    .A2(_06502_),
    .B1(_06984_),
    .X(_06985_));
 sky130_fd_sc_hd__a2bb2oi_1 _12841_ (.A1_N(_06955_),
    .A2_N(_06985_),
    .B1(_06955_),
    .B2(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__buf_1 _12842_ (.A(\e1.alu1.a[5] ),
    .X(_06987_));
 sky130_fd_sc_hd__buf_1 _12843_ (.A(_06495_),
    .X(_06988_));
 sky130_fd_sc_hd__o21a_1 _12844_ (.A1(_00039_),
    .A2(_06988_),
    .B1(_06570_),
    .X(_06989_));
 sky130_fd_sc_hd__o22ai_1 _12845_ (.A1(_06987_),
    .A2(_06494_),
    .B1(_06719_),
    .B2(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__or2_1 _12846_ (.A(_00275_),
    .B(_06682_),
    .X(_00200_));
 sky130_fd_sc_hd__or3_1 _12847_ (.A(_00039_),
    .B(_06988_),
    .C(_06945_),
    .X(_06991_));
 sky130_fd_sc_hd__o221a_1 _12848_ (.A1(_00195_),
    .A2(_06943_),
    .B1(_06966_),
    .B2(_00200_),
    .C1(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__o211ai_1 _12849_ (.A1(_06587_),
    .A2(_06986_),
    .B1(_06990_),
    .C1(_06992_),
    .Y(_00201_));
 sky130_fd_sc_hd__or2_1 _12850_ (.A(_00266_),
    .B(_06972_),
    .X(_06993_));
 sky130_fd_sc_hd__clkbuf_2 _12851_ (.A(_06993_),
    .X(_00187_));
 sky130_fd_sc_hd__buf_1 _12852_ (.A(_06501_),
    .X(_06994_));
 sky130_fd_sc_hd__o32a_1 _12853_ (.A1(_06994_),
    .A2(_00038_),
    .A3(_06949_),
    .B1(_00182_),
    .B2(_06975_),
    .X(_06995_));
 sky130_fd_sc_hd__clkbuf_2 _12854_ (.A(_06503_),
    .X(_06996_));
 sky130_fd_sc_hd__o21a_1 _12855_ (.A1(_06994_),
    .A2(_00038_),
    .B1(_06979_),
    .X(_06997_));
 sky130_fd_sc_hd__o22ai_4 _12856_ (.A1(_06558_),
    .A2(_06996_),
    .B1(_06978_),
    .B2(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__o211ai_4 _12857_ (.A1(_06957_),
    .A2(_06956_),
    .B1(_06655_),
    .C1(_06984_),
    .Y(_06999_));
 sky130_fd_sc_hd__o2111ai_4 _12858_ (.A1(_06971_),
    .A2(_00187_),
    .B1(_06995_),
    .C1(_06998_),
    .D1(_06999_),
    .Y(_00188_));
 sky130_fd_sc_hd__inv_2 _12859_ (.A(_00197_),
    .Y(_00198_));
 sky130_fd_sc_hd__or2_1 _12860_ (.A(_06705_),
    .B(_00257_),
    .X(_07000_));
 sky130_fd_sc_hd__buf_1 _12861_ (.A(_07000_),
    .X(_00174_));
 sky130_fd_sc_hd__buf_2 _12862_ (.A(_06460_),
    .X(_00034_));
 sky130_fd_sc_hd__inv_2 _12863_ (.A(_06464_),
    .Y(_07001_));
 sky130_fd_sc_hd__o22a_1 _12864_ (.A1(_00034_),
    .A2(_06462_),
    .B1(_06470_),
    .B2(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__a2bb2oi_2 _12865_ (.A1_N(_06459_),
    .A2_N(_07002_),
    .B1(_06459_),
    .B2(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__buf_1 _12866_ (.A(\e1.alu1.a[3] ),
    .X(_07004_));
 sky130_fd_sc_hd__nor2_1 _12867_ (.A(_06455_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__a21oi_2 _12868_ (.A1(_06563_),
    .A2(_07004_),
    .B1(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__inv_2 _12869_ (.A(_07006_),
    .Y(_07007_));
 sky130_fd_sc_hd__o32a_1 _12870_ (.A1(_06456_),
    .A2(_00035_),
    .A3(_06576_),
    .B1(_00171_),
    .B2(_06912_),
    .X(_07008_));
 sky130_fd_sc_hd__o221a_1 _12871_ (.A1(_06852_),
    .A2(_07007_),
    .B1(_06675_),
    .B2(_07005_),
    .C1(_07008_),
    .X(_07009_));
 sky130_fd_sc_hd__o221ai_4 _12872_ (.A1(_06884_),
    .A2(_00174_),
    .B1(_06845_),
    .B2(_07003_),
    .C1(_07009_),
    .Y(_00175_));
 sky130_fd_sc_hd__inv_2 _12873_ (.A(_00184_),
    .Y(_00185_));
 sky130_fd_sc_hd__nor2_2 _12874_ (.A(_06653_),
    .B(_06472_),
    .Y(_07010_));
 sky130_fd_sc_hd__nor2_2 _12875_ (.A(_06461_),
    .B(_00034_),
    .Y(_07011_));
 sky130_fd_sc_hd__o21a_1 _12876_ (.A1(_06852_),
    .A2(_07011_),
    .B1(_06619_),
    .X(_07012_));
 sky130_fd_sc_hd__a22o_1 _12877_ (.A1(_06471_),
    .A2(_06464_),
    .B1(_06470_),
    .B2(_07001_),
    .X(_07013_));
 sky130_fd_sc_hd__or2_1 _12878_ (.A(_06565_),
    .B(_00248_),
    .X(_00155_));
 sky130_fd_sc_hd__nand2_1 _12879_ (.A(_06910_),
    .B(_07011_),
    .Y(_07014_));
 sky130_fd_sc_hd__o221a_1 _12880_ (.A1(_00151_),
    .A2(_06912_),
    .B1(_06944_),
    .B2(_00155_),
    .C1(_07014_),
    .X(_07015_));
 sky130_fd_sc_hd__o221ai_2 _12881_ (.A1(_07010_),
    .A2(_07012_),
    .B1(_06845_),
    .B2(_07013_),
    .C1(_07015_),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_2 _12882_ (.A(_00152_),
    .Y(_00153_));
 sky130_fd_sc_hd__or2_1 _12883_ (.A(_06972_),
    .B(_00239_),
    .X(_07016_));
 sky130_fd_sc_hd__buf_1 _12884_ (.A(_07016_),
    .X(_00133_));
 sky130_fd_sc_hd__clkbuf_4 _12885_ (.A(_06466_),
    .X(_00032_));
 sky130_fd_sc_hd__buf_1 _12886_ (.A(_06969_),
    .X(_07017_));
 sky130_fd_sc_hd__o32a_1 _12887_ (.A1(_07017_),
    .A2(_00032_),
    .A3(_06602_),
    .B1(_00130_),
    .B2(_06975_),
    .X(_07018_));
 sky130_fd_sc_hd__clkbuf_2 _12888_ (.A(\e1.alu1.a[1] ),
    .X(_07019_));
 sky130_fd_sc_hd__o21a_1 _12889_ (.A1(_07017_),
    .A2(_00032_),
    .B1(_06979_),
    .X(_07020_));
 sky130_fd_sc_hd__o22ai_4 _12890_ (.A1(_06708_),
    .A2(_07019_),
    .B1(_06978_),
    .B2(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__inv_2 _12891_ (.A(_00135_),
    .Y(_07022_));
 sky130_fd_sc_hd__inv_2 _12892_ (.A(_06469_),
    .Y(_07023_));
 sky130_fd_sc_hd__a221o_1 _12893_ (.A1(_07022_),
    .A2(_07023_),
    .B1(_00135_),
    .B2(_06469_),
    .C1(_06862_),
    .X(_07024_));
 sky130_fd_sc_hd__o2111ai_4 _12894_ (.A1(_06971_),
    .A2(_00133_),
    .B1(_07018_),
    .C1(_07021_),
    .D1(_07024_),
    .Y(_00136_));
 sky130_fd_sc_hd__o22a_1 _12895_ (.A1(_06716_),
    .A2(\e1.alu1.a[30] ),
    .B1(_06712_),
    .B2(_06709_),
    .X(_07025_));
 sky130_fd_sc_hd__or2_2 _12896_ (.A(_06743_),
    .B(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__o22a_1 _12897_ (.A1(_06687_),
    .A2(_06694_),
    .B1(_06688_),
    .B2(_06685_),
    .X(_07027_));
 sky130_fd_sc_hd__o21bai_1 _12898_ (.A1(_06671_),
    .A2(_06674_),
    .B1_N(_07027_),
    .Y(_07028_));
 sky130_fd_sc_hd__o32a_1 _12899_ (.A1(_06270_),
    .A2(_06571_),
    .A3(_06609_),
    .B1(_06600_),
    .B2(_06597_),
    .X(_07029_));
 sky130_fd_sc_hd__o22a_1 _12900_ (.A1(_06621_),
    .A2(_06613_),
    .B1(_06615_),
    .B2(_07029_),
    .X(_07030_));
 sky130_fd_sc_hd__o22a_1 _12901_ (.A1(_06646_),
    .A2(_06644_),
    .B1(_06650_),
    .B2(_07030_),
    .X(_07031_));
 sky130_fd_sc_hd__or3_1 _12902_ (.A(_06663_),
    .B(_06666_),
    .C(_07027_),
    .X(_07032_));
 sky130_fd_sc_hd__o221a_1 _12903_ (.A1(_06697_),
    .A2(_06694_),
    .B1(_07028_),
    .B2(_07031_),
    .C1(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__or4_4 _12904_ (.A(_06572_),
    .B(_06615_),
    .C(_06609_),
    .D(_06650_),
    .X(_07034_));
 sky130_fd_sc_hd__or3_4 _12905_ (.A(_07026_),
    .B(_07028_),
    .C(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__or2_1 _12906_ (.A(_06810_),
    .B(_06816_),
    .X(_07036_));
 sky130_fd_sc_hd__o22a_1 _12907_ (.A1(_06377_),
    .A2(\e1.alu1.a1.b[16] ),
    .B1(_06371_),
    .B2(_06856_),
    .X(_07037_));
 sky130_fd_sc_hd__or4_4 _12908_ (.A(_06832_),
    .B(_06853_),
    .C(_06787_),
    .D(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__or4_4 _12909_ (.A(_06795_),
    .B(_06839_),
    .C(_07036_),
    .D(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__o22a_1 _12910_ (.A1(_06872_),
    .A2(_06390_),
    .B1(_06523_),
    .B2(_06391_),
    .X(_07040_));
 sky130_fd_sc_hd__o22a_1 _12911_ (.A1(_06399_),
    .A2(_06889_),
    .B1(_06402_),
    .B2(_06398_),
    .X(_07041_));
 sky130_fd_sc_hd__o22a_1 _12912_ (.A1(_06899_),
    .A2(_06416_),
    .B1(_06415_),
    .B2(_06417_),
    .X(_07042_));
 sky130_fd_sc_hd__or2_1 _12913_ (.A(_06907_),
    .B(_06908_),
    .X(_07043_));
 sky130_fd_sc_hd__or4b_4 _12914_ (.A(_07040_),
    .B(_07041_),
    .C(_07042_),
    .D_N(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__o22a_1 _12915_ (.A1(_06939_),
    .A2(_06448_),
    .B1(_06447_),
    .B2(_06449_),
    .X(_07045_));
 sky130_fd_sc_hd__o22a_1 _12916_ (.A1(_06922_),
    .A2(_06423_),
    .B1(_06517_),
    .B2(_06424_),
    .X(_07046_));
 sky130_fd_sc_hd__o22a_1 _12917_ (.A1(_06951_),
    .A2(_06439_),
    .B1(_06936_),
    .B2(_06948_),
    .X(_07047_));
 sky130_fd_sc_hd__o22a_1 _12918_ (.A1(_06931_),
    .A2(_06431_),
    .B1(_06430_),
    .B2(_06432_),
    .X(_07048_));
 sky130_fd_sc_hd__or4_4 _12919_ (.A(_07045_),
    .B(_07046_),
    .C(_07047_),
    .D(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__o22a_1 _12920_ (.A1(_06987_),
    .A2(_06494_),
    .B1(_06492_),
    .B2(_06495_),
    .X(_07050_));
 sky130_fd_sc_hd__o22a_1 _12921_ (.A1(_06500_),
    .A2(_06996_),
    .B1(_06994_),
    .B2(_06983_),
    .X(_07051_));
 sky130_fd_sc_hd__o22a_1 _12922_ (.A1(_06977_),
    .A2(_06486_),
    .B1(_06485_),
    .B2(_06487_),
    .X(_07052_));
 sky130_fd_sc_hd__o22a_1 _12923_ (.A1(_06962_),
    .A2(_06478_),
    .B1(_06477_),
    .B2(_06479_),
    .X(_07053_));
 sky130_fd_sc_hd__or4_4 _12924_ (.A(_07050_),
    .B(_07051_),
    .C(_07052_),
    .D(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__o21ai_1 _12925_ (.A1(_07010_),
    .A2(_07011_),
    .B1(_07007_),
    .Y(_07055_));
 sky130_fd_sc_hd__or2_1 _12926_ (.A(_06969_),
    .B(_00024_),
    .X(_07056_));
 sky130_fd_sc_hd__inv_2 _12927_ (.A(_06970_),
    .Y(_00094_));
 sky130_fd_sc_hd__a21o_1 _12928_ (.A1(_07019_),
    .A2(_07056_),
    .B1(_00094_),
    .X(_07057_));
 sky130_fd_sc_hd__or3_2 _12929_ (.A(_06935_),
    .B(_06472_),
    .C(_07006_),
    .X(_07058_));
 sky130_fd_sc_hd__o221a_1 _12930_ (.A1(_06456_),
    .A2(_07004_),
    .B1(_07055_),
    .B2(_07057_),
    .C1(_07058_),
    .X(_07059_));
 sky130_fd_sc_hd__o32a_1 _12931_ (.A1(_06501_),
    .A2(_06996_),
    .A3(_07050_),
    .B1(_06987_),
    .B2(_06988_),
    .X(_07060_));
 sky130_fd_sc_hd__o22a_1 _12932_ (.A1(_06977_),
    .A2(_06974_),
    .B1(_07052_),
    .B2(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__or2_1 _12933_ (.A(_07053_),
    .B(_07061_),
    .X(_07062_));
 sky130_fd_sc_hd__o221a_1 _12934_ (.A1(_07054_),
    .A2(_07059_),
    .B1(_06962_),
    .B2(_06963_),
    .C1(_07062_),
    .X(_07063_));
 sky130_fd_sc_hd__o32a_1 _12935_ (.A1(_06951_),
    .A2(_06440_),
    .A3(_07045_),
    .B1(_06939_),
    .B2(_06940_),
    .X(_07064_));
 sky130_fd_sc_hd__o22a_1 _12936_ (.A1(_06931_),
    .A2(_06929_),
    .B1(_07048_),
    .B2(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__or2_1 _12937_ (.A(_07046_),
    .B(_07065_),
    .X(_07066_));
 sky130_fd_sc_hd__o221a_1 _12938_ (.A1(_06922_),
    .A2(_06924_),
    .B1(_07049_),
    .B2(_07063_),
    .C1(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__o32a_1 _12939_ (.A1(_06411_),
    .A2(_06409_),
    .A3(_07042_),
    .B1(_06899_),
    .B2(_06900_),
    .X(_07068_));
 sky130_fd_sc_hd__o22a_1 _12940_ (.A1(_06886_),
    .A2(_06889_),
    .B1(_07041_),
    .B2(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__or2_1 _12941_ (.A(_07040_),
    .B(_07069_),
    .X(_07070_));
 sky130_fd_sc_hd__o221a_1 _12942_ (.A1(_06872_),
    .A2(_06873_),
    .B1(_07044_),
    .B2(_07067_),
    .C1(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__o32a_1 _12943_ (.A1(_06377_),
    .A2(_06856_),
    .A3(_06853_),
    .B1(_06848_),
    .B2(_06850_),
    .X(_07072_));
 sky130_fd_sc_hd__o22a_1 _12944_ (.A1(_06836_),
    .A2(_06838_),
    .B1(_06839_),
    .B2(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__o22a_1 _12945_ (.A1(_06828_),
    .A2(_06830_),
    .B1(_06832_),
    .B2(_07073_),
    .X(_07074_));
 sky130_fd_sc_hd__or3_1 _12946_ (.A(_06814_),
    .B(_06815_),
    .C(_06810_),
    .X(_07075_));
 sky130_fd_sc_hd__o221a_1 _12947_ (.A1(_06804_),
    .A2(_06807_),
    .B1(_07036_),
    .B2(_07074_),
    .C1(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__o22a_1 _12948_ (.A1(_06791_),
    .A2(_06794_),
    .B1(_06795_),
    .B2(_07076_),
    .X(_07077_));
 sky130_fd_sc_hd__or2_1 _12949_ (.A(_06787_),
    .B(_07077_),
    .X(_07078_));
 sky130_fd_sc_hd__o221a_1 _12950_ (.A1(_06782_),
    .A2(_06784_),
    .B1(_07039_),
    .B2(_07071_),
    .C1(_07078_),
    .X(_07079_));
 sky130_fd_sc_hd__or3_4 _12951_ (.A(_06713_),
    .B(_06717_),
    .C(_06743_),
    .X(_07080_));
 sky130_fd_sc_hd__o221ai_4 _12952_ (.A1(_07026_),
    .A2(_07033_),
    .B1(_07035_),
    .B2(_07079_),
    .C1(_07080_),
    .Y(_07081_));
 sky130_fd_sc_hd__o22a_1 _12953_ (.A1(_06707_),
    .A2(_07019_),
    .B1(_07017_),
    .B2(_06466_),
    .X(_07082_));
 sky130_fd_sc_hd__buf_1 _12954_ (.A(\e1.alu1.a[0] ),
    .X(_07083_));
 sky130_fd_sc_hd__nand2_1 _12955_ (.A(\e1.alu1.a1.b[0] ),
    .B(_07083_),
    .Y(_07084_));
 sky130_fd_sc_hd__o21a_1 _12956_ (.A1(_06734_),
    .A2(_07083_),
    .B1(_07084_),
    .X(_07085_));
 sky130_fd_sc_hd__or4_4 _12957_ (.A(_07082_),
    .B(_07085_),
    .C(_07055_),
    .D(_07044_),
    .X(_07086_));
 sky130_fd_sc_hd__or2_1 _12958_ (.A(_07049_),
    .B(_07054_),
    .X(_07087_));
 sky130_fd_sc_hd__or4_4 _12959_ (.A(_07086_),
    .B(_07087_),
    .C(_07035_),
    .D(_07039_),
    .X(_07088_));
 sky130_fd_sc_hd__o221a_2 _12960_ (.A1(_06744_),
    .A2(_07081_),
    .B1(_06735_),
    .B2(_06738_),
    .C1(_07088_),
    .X(_00027_));
 sky130_fd_sc_hd__inv_2 _12961_ (.A(_00027_),
    .Y(_07089_));
 sky130_fd_sc_hd__nor2_2 _12962_ (.A(_06736_),
    .B(_06738_),
    .Y(_07090_));
 sky130_fd_sc_hd__buf_2 _12963_ (.A(_07088_),
    .X(_00021_));
 sky130_fd_sc_hd__o21ai_4 _12964_ (.A1(_07090_),
    .A2(_07081_),
    .B1(_00021_),
    .Y(_07091_));
 sky130_fd_sc_hd__o21a_1 _12965_ (.A1(_06654_),
    .A2(_06891_),
    .B1(_07084_),
    .X(_07092_));
 sky130_fd_sc_hd__o22ai_1 _12966_ (.A1(_06734_),
    .A2(_07083_),
    .B1(_06695_),
    .B2(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__or2_1 _12967_ (.A(_06583_),
    .B(_00230_),
    .X(_00095_));
 sky130_fd_sc_hd__o32a_1 _12968_ (.A1(_00030_),
    .A2(_06276_),
    .A3(_03680_),
    .B1(_00093_),
    .B2(_06911_),
    .X(_07094_));
 sky130_fd_sc_hd__o221a_1 _12969_ (.A1(_06792_),
    .A2(_07084_),
    .B1(_06879_),
    .B2(_00095_),
    .C1(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__o311a_1 _12970_ (.A1(_06566_),
    .A2(_06578_),
    .A3(_07091_),
    .B1(_07093_),
    .C1(_07095_),
    .X(_07096_));
 sky130_fd_sc_hd__o31ai_1 _12971_ (.A1(_06578_),
    .A2(_06303_),
    .A3(_07089_),
    .B1(_07096_),
    .Y(_00099_));
 sky130_fd_sc_hd__inv_2 _12972_ (.A(_07091_),
    .Y(_00025_));
 sky130_fd_sc_hd__and3_1 _12973_ (.A(_06297_),
    .B(_06282_),
    .C(_06299_),
    .X(_00023_));
 sky130_fd_sc_hd__or3b_1 _12974_ (.A(_00023_),
    .B(_06276_),
    .C_N(_00096_),
    .X(_00097_));
 sky130_fd_sc_hd__inv_2 _12975_ (.A(_06283_),
    .Y(_07097_));
 sky130_fd_sc_hd__a311oi_4 _12976_ (.A1(_03966_),
    .A2(_07097_),
    .A3(_00021_),
    .B1(_00028_),
    .C1(_00026_),
    .Y(_00029_));
 sky130_fd_sc_hd__clkbuf_1 _12977_ (.A(_06297_),
    .X(_07098_));
 sky130_fd_sc_hd__nor2_1 _12978_ (.A(_07098_),
    .B(_07097_),
    .Y(_00022_));
 sky130_fd_sc_hd__nor2_8 _12979_ (.A(_06551_),
    .B(_06290_),
    .Y(_00020_));
 sky130_fd_sc_hd__and3_1 _12980_ (.A(_07098_),
    .B(_03969_),
    .C(_03971_),
    .X(_00016_));
 sky130_fd_sc_hd__a21o_1 _12981_ (.A1(_00004_),
    .A2(_06299_),
    .B1(_00016_),
    .X(_00017_));
 sky130_fd_sc_hd__inv_2 _12982_ (.A(_06284_),
    .Y(_00009_));
 sky130_fd_sc_hd__nor3_4 _12983_ (.A(\c1.instruction2[29] ),
    .B(\c1.instruction2[30] ),
    .C(_06287_),
    .Y(_00012_));
 sky130_fd_sc_hd__and3_1 _12984_ (.A(_07098_),
    .B(_06282_),
    .C(_03971_),
    .X(_00008_));
 sky130_fd_sc_hd__inv_2 _12985_ (.A(_03500_),
    .Y(_07099_));
 sky130_fd_sc_hd__nor2_1 _12986_ (.A(_03927_),
    .B(_07099_),
    .Y(_00003_));
 sky130_fd_sc_hd__o22a_1 _12987_ (.A1(_03934_),
    .A2(\c1.instruction1[22] ),
    .B1(\c1.instruction2[9] ),
    .B2(_00400_),
    .X(_07100_));
 sky130_fd_sc_hd__o221a_1 _12988_ (.A1(\c1.instruction2[11] ),
    .A2(_00406_),
    .B1(_03929_),
    .B2(net50),
    .C1(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__o22a_1 _12989_ (.A1(\c1.instruction2[7] ),
    .A2(_03858_),
    .B1(\c1.instruction2[10] ),
    .B2(_03842_),
    .X(_07102_));
 sky130_fd_sc_hd__o221a_1 _12990_ (.A1(_03928_),
    .A2(net53),
    .B1(_03931_),
    .B2(net40),
    .C1(_07102_),
    .X(_07103_));
 sky130_fd_sc_hd__o221a_1 _12991_ (.A1(\c1.instruction2[8] ),
    .A2(_00397_),
    .B1(_03935_),
    .B2(\c1.instruction1[23] ),
    .C1(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__a21oi_1 _12992_ (.A1(_07101_),
    .A2(_07104_),
    .B1(_07099_),
    .Y(_00002_));
 sky130_fd_sc_hd__nor2_1 _12993_ (.A(_03938_),
    .B(_07099_),
    .Y(_00001_));
 sky130_fd_sc_hd__clkbuf_1 _12994_ (.A(_03500_),
    .X(_00000_));
 sky130_fd_sc_hd__inv_2 _12995_ (.A(\e1.pc[0] ),
    .Y(_01210_));
 sky130_fd_sc_hd__inv_2 _12996_ (.A(\e1.pc[1] ),
    .Y(_01212_));
 sky130_fd_sc_hd__inv_2 _12997_ (.A(\e1.pc[2] ),
    .Y(_01214_));
 sky130_fd_sc_hd__inv_2 _12998_ (.A(\e1.pc[3] ),
    .Y(_01216_));
 sky130_fd_sc_hd__inv_2 _12999_ (.A(\e1.pc[4] ),
    .Y(_01218_));
 sky130_fd_sc_hd__inv_2 _13000_ (.A(\e1.pc[5] ),
    .Y(_01220_));
 sky130_fd_sc_hd__inv_2 _13001_ (.A(\e1.pc[6] ),
    .Y(_01222_));
 sky130_fd_sc_hd__inv_2 _13002_ (.A(\e1.pc[7] ),
    .Y(_01224_));
 sky130_fd_sc_hd__inv_2 _13003_ (.A(\e1.pc[8] ),
    .Y(_01226_));
 sky130_fd_sc_hd__inv_2 _13004_ (.A(\e1.pc[9] ),
    .Y(_01228_));
 sky130_fd_sc_hd__inv_2 _13005_ (.A(\e1.pc[10] ),
    .Y(_01230_));
 sky130_fd_sc_hd__inv_2 _13006_ (.A(\e1.pc[11] ),
    .Y(_01232_));
 sky130_fd_sc_hd__inv_2 _13007_ (.A(\e1.pc[12] ),
    .Y(_01234_));
 sky130_fd_sc_hd__inv_2 _13008_ (.A(\e1.pc[13] ),
    .Y(_01236_));
 sky130_fd_sc_hd__inv_2 _13009_ (.A(\e1.pc[14] ),
    .Y(_01238_));
 sky130_fd_sc_hd__inv_2 _13010_ (.A(\e1.pc[15] ),
    .Y(_01240_));
 sky130_fd_sc_hd__inv_2 _13011_ (.A(\e1.pc[16] ),
    .Y(_01242_));
 sky130_fd_sc_hd__inv_2 _13012_ (.A(\e1.pc[17] ),
    .Y(_01244_));
 sky130_fd_sc_hd__inv_2 _13013_ (.A(\e1.pc[18] ),
    .Y(_01246_));
 sky130_fd_sc_hd__inv_2 _13014_ (.A(\e1.pc[19] ),
    .Y(_01248_));
 sky130_fd_sc_hd__inv_2 _13015_ (.A(\e1.pc[20] ),
    .Y(_01250_));
 sky130_fd_sc_hd__inv_2 _13016_ (.A(\e1.pc[21] ),
    .Y(_01252_));
 sky130_fd_sc_hd__inv_2 _13017_ (.A(\e1.pc[22] ),
    .Y(_01254_));
 sky130_fd_sc_hd__inv_2 _13018_ (.A(\e1.pc[23] ),
    .Y(_01256_));
 sky130_fd_sc_hd__inv_2 _13019_ (.A(\e1.pc[24] ),
    .Y(_01258_));
 sky130_fd_sc_hd__inv_2 _13020_ (.A(\e1.pc[25] ),
    .Y(_01260_));
 sky130_fd_sc_hd__inv_2 _13021_ (.A(\e1.pc[26] ),
    .Y(_01262_));
 sky130_fd_sc_hd__inv_2 _13022_ (.A(\e1.pc[27] ),
    .Y(_01264_));
 sky130_fd_sc_hd__inv_2 _13023_ (.A(\e1.pc[28] ),
    .Y(_01266_));
 sky130_fd_sc_hd__inv_2 _13024_ (.A(\e1.pc[29] ),
    .Y(_01268_));
 sky130_fd_sc_hd__inv_2 _13025_ (.A(\e1.pc[30] ),
    .Y(_01270_));
 sky130_fd_sc_hd__o221a_1 _13026_ (.A1(\next_pc[1] ),
    .A2(_03665_),
    .B1(_06756_),
    .B2(_03669_),
    .C1(_03740_),
    .X(_03663_));
 sky130_fd_sc_hd__mux2_1 _13027_ (.A0(wdata[0]),
    .A1(rdata[0]),
    .S(net7),
    .X(\wbmemout[0] ));
 sky130_fd_sc_hd__mux2_1 _13028_ (.A0(wdata[1]),
    .A1(rdata[1]),
    .S(net7),
    .X(\wbmemout[1] ));
 sky130_fd_sc_hd__mux2_1 _13029_ (.A0(wdata[2]),
    .A1(rdata[2]),
    .S(net7),
    .X(\wbmemout[2] ));
 sky130_fd_sc_hd__mux2_1 _13030_ (.A0(wdata[3]),
    .A1(rdata[3]),
    .S(net7),
    .X(\wbmemout[3] ));
 sky130_fd_sc_hd__mux2_1 _13031_ (.A0(wdata[4]),
    .A1(rdata[4]),
    .S(net7),
    .X(\wbmemout[4] ));
 sky130_fd_sc_hd__mux2_4 _13032_ (.A0(wdata[5]),
    .A1(rdata[5]),
    .S(net7),
    .X(\wbmemout[5] ));
 sky130_fd_sc_hd__mux2_1 _13033_ (.A0(wdata[6]),
    .A1(rdata[6]),
    .S(net7),
    .X(\wbmemout[6] ));
 sky130_fd_sc_hd__mux2_1 _13034_ (.A0(wdata[7]),
    .A1(rdata[7]),
    .S(net7),
    .X(\wbmemout[7] ));
 sky130_fd_sc_hd__mux2_4 _13035_ (.A0(wdata[8]),
    .A1(rdata[8]),
    .S(net7),
    .X(\wbmemout[8] ));
 sky130_fd_sc_hd__mux2_2 _13036_ (.A0(wdata[9]),
    .A1(rdata[9]),
    .S(net6),
    .X(\wbmemout[9] ));
 sky130_fd_sc_hd__mux2_4 _13037_ (.A0(wdata[10]),
    .A1(rdata[10]),
    .S(ren),
    .X(\wbmemout[10] ));
 sky130_fd_sc_hd__mux2_2 _13038_ (.A0(wdata[11]),
    .A1(rdata[11]),
    .S(ren),
    .X(\wbmemout[11] ));
 sky130_fd_sc_hd__mux2_1 _13039_ (.A0(wdata[12]),
    .A1(rdata[12]),
    .S(ren),
    .X(\wbmemout[12] ));
 sky130_fd_sc_hd__mux2_1 _13040_ (.A0(wdata[13]),
    .A1(rdata[13]),
    .S(ren),
    .X(\wbmemout[13] ));
 sky130_fd_sc_hd__mux2_1 _13041_ (.A0(wdata[14]),
    .A1(rdata[14]),
    .S(ren),
    .X(\wbmemout[14] ));
 sky130_fd_sc_hd__mux2_1 _13042_ (.A0(wdata[15]),
    .A1(rdata[15]),
    .S(ren),
    .X(\wbmemout[15] ));
 sky130_fd_sc_hd__mux2_1 _13043_ (.A0(wdata[16]),
    .A1(rdata[16]),
    .S(ren),
    .X(\wbmemout[16] ));
 sky130_fd_sc_hd__mux2_1 _13044_ (.A0(wdata[17]),
    .A1(rdata[17]),
    .S(ren),
    .X(\wbmemout[17] ));
 sky130_fd_sc_hd__mux2_1 _13045_ (.A0(wdata[18]),
    .A1(rdata[18]),
    .S(net7),
    .X(\wbmemout[18] ));
 sky130_fd_sc_hd__mux2_1 _13046_ (.A0(wdata[19]),
    .A1(rdata[19]),
    .S(net7),
    .X(\wbmemout[19] ));
 sky130_fd_sc_hd__mux2_1 _13047_ (.A0(wdata[20]),
    .A1(rdata[20]),
    .S(net6),
    .X(\wbmemout[20] ));
 sky130_fd_sc_hd__mux2_1 _13048_ (.A0(wdata[21]),
    .A1(rdata[21]),
    .S(net6),
    .X(\wbmemout[21] ));
 sky130_fd_sc_hd__mux2_1 _13049_ (.A0(wdata[22]),
    .A1(rdata[22]),
    .S(net6),
    .X(\wbmemout[22] ));
 sky130_fd_sc_hd__mux2_1 _13050_ (.A0(wdata[23]),
    .A1(rdata[23]),
    .S(net6),
    .X(\wbmemout[23] ));
 sky130_fd_sc_hd__mux2_1 _13051_ (.A0(wdata[24]),
    .A1(rdata[24]),
    .S(net6),
    .X(\wbmemout[24] ));
 sky130_fd_sc_hd__mux2_1 _13052_ (.A0(wdata[25]),
    .A1(rdata[25]),
    .S(net6),
    .X(\wbmemout[25] ));
 sky130_fd_sc_hd__mux2_1 _13053_ (.A0(wdata[26]),
    .A1(rdata[26]),
    .S(net6),
    .X(\wbmemout[26] ));
 sky130_fd_sc_hd__mux2_1 _13054_ (.A0(wdata[27]),
    .A1(rdata[27]),
    .S(net6),
    .X(\wbmemout[27] ));
 sky130_fd_sc_hd__mux2_1 _13055_ (.A0(wdata[28]),
    .A1(rdata[28]),
    .S(net6),
    .X(\wbmemout[28] ));
 sky130_fd_sc_hd__mux2_1 _13056_ (.A0(wdata[29]),
    .A1(rdata[29]),
    .S(net6),
    .X(\wbmemout[29] ));
 sky130_fd_sc_hd__mux2_1 _13057_ (.A0(wdata[30]),
    .A1(rdata[30]),
    .S(net6),
    .X(\wbmemout[30] ));
 sky130_fd_sc_hd__mux2_1 _13058_ (.A0(wdata[31]),
    .A1(rdata[31]),
    .S(net7),
    .X(\wbmemout[31] ));
 sky130_fd_sc_hd__mux2_4 _13059_ (.A0(_00099_),
    .A1(\e1.alu1.a1.b[0] ),
    .S(_00020_),
    .X(\e1.alu1.out[0] ));
 sky130_fd_sc_hd__mux2_1 _13060_ (.A0(_00136_),
    .A1(\e1.alu1.a1.b[1] ),
    .S(_00020_),
    .X(\e1.alu1.out[1] ));
 sky130_fd_sc_hd__mux2_2 _13061_ (.A0(_00156_),
    .A1(\e1.alu1.a1.b[2] ),
    .S(_00020_),
    .X(\e1.alu1.out[2] ));
 sky130_fd_sc_hd__mux2_1 _13062_ (.A0(_00175_),
    .A1(\e1.alu1.a1.b[3] ),
    .S(net1),
    .X(\e1.alu1.out[3] ));
 sky130_fd_sc_hd__mux2_2 _13063_ (.A0(_00188_),
    .A1(\e1.alu1.a1.b[4] ),
    .S(net1),
    .X(\e1.alu1.out[4] ));
 sky130_fd_sc_hd__mux2_1 _13064_ (.A0(_00201_),
    .A1(\e1.alu1.a1.b[5] ),
    .S(net1),
    .X(\e1.alu1.out[5] ));
 sky130_fd_sc_hd__mux2_2 _13065_ (.A0(_00214_),
    .A1(\e1.alu1.a1.b[6] ),
    .S(_00020_),
    .X(\e1.alu1.out[6] ));
 sky130_fd_sc_hd__mux2_2 _13066_ (.A0(_00226_),
    .A1(\e1.alu1.a1.b[7] ),
    .S(_00020_),
    .X(\e1.alu1.out[7] ));
 sky130_fd_sc_hd__mux2_2 _13067_ (.A0(_00235_),
    .A1(\e1.alu1.a1.b[8] ),
    .S(_00020_),
    .X(\e1.alu1.out[8] ));
 sky130_fd_sc_hd__mux2_1 _13068_ (.A0(_00244_),
    .A1(\e1.alu1.a1.b[9] ),
    .S(_00020_),
    .X(\e1.alu1.out[9] ));
 sky130_fd_sc_hd__mux2_1 _13069_ (.A0(_00253_),
    .A1(\e1.alu1.a1.b[10] ),
    .S(_00020_),
    .X(\e1.alu1.out[10] ));
 sky130_fd_sc_hd__mux2_1 _13070_ (.A0(_00262_),
    .A1(\e1.alu1.a1.b[11] ),
    .S(_00020_),
    .X(\e1.alu1.out[11] ));
 sky130_fd_sc_hd__mux2_1 _13071_ (.A0(_00271_),
    .A1(\e1.alu1.a1.b[12] ),
    .S(_00020_),
    .X(\e1.alu1.out[12] ));
 sky130_fd_sc_hd__mux2_1 _13072_ (.A0(_00280_),
    .A1(\e1.alu1.a1.b[13] ),
    .S(_00020_),
    .X(\e1.alu1.out[13] ));
 sky130_fd_sc_hd__mux2_1 _13073_ (.A0(_00289_),
    .A1(\e1.alu1.a1.b[14] ),
    .S(_00020_),
    .X(\e1.alu1.out[14] ));
 sky130_fd_sc_hd__mux2_1 _13074_ (.A0(_00297_),
    .A1(\e1.alu1.a1.b[15] ),
    .S(_00020_),
    .X(\e1.alu1.out[15] ));
 sky130_fd_sc_hd__mux2_1 _13075_ (.A0(_00303_),
    .A1(\e1.alu1.a1.b[16] ),
    .S(_00020_),
    .X(\e1.alu1.out[16] ));
 sky130_fd_sc_hd__mux2_2 _13076_ (.A0(_00309_),
    .A1(\e1.alu1.a1.b[17] ),
    .S(_00020_),
    .X(\e1.alu1.out[17] ));
 sky130_fd_sc_hd__mux2_1 _13077_ (.A0(_00315_),
    .A1(\e1.alu1.a1.b[18] ),
    .S(net1),
    .X(\e1.alu1.out[18] ));
 sky130_fd_sc_hd__mux2_1 _13078_ (.A0(_00321_),
    .A1(\e1.alu1.a1.b[19] ),
    .S(net1),
    .X(\e1.alu1.out[19] ));
 sky130_fd_sc_hd__mux2_1 _13079_ (.A0(_00327_),
    .A1(\e1.alu1.a1.b[20] ),
    .S(net1),
    .X(\e1.alu1.out[20] ));
 sky130_fd_sc_hd__mux2_1 _13080_ (.A0(_00333_),
    .A1(\e1.alu1.a1.b[21] ),
    .S(net1),
    .X(\e1.alu1.out[21] ));
 sky130_fd_sc_hd__mux2_1 _13081_ (.A0(_00339_),
    .A1(\e1.alu1.a1.b[22] ),
    .S(net1),
    .X(\e1.alu1.out[22] ));
 sky130_fd_sc_hd__mux2_1 _13082_ (.A0(_00345_),
    .A1(\e1.alu1.a1.b[23] ),
    .S(net1),
    .X(\e1.alu1.out[23] ));
 sky130_fd_sc_hd__mux2_1 _13083_ (.A0(_00351_),
    .A1(\e1.alu1.a1.b[24] ),
    .S(net1),
    .X(\e1.alu1.out[24] ));
 sky130_fd_sc_hd__mux2_1 _13084_ (.A0(_00357_),
    .A1(\e1.alu1.a1.b[25] ),
    .S(net1),
    .X(\e1.alu1.out[25] ));
 sky130_fd_sc_hd__mux2_1 _13085_ (.A0(_00363_),
    .A1(\e1.alu1.a1.b[26] ),
    .S(net1),
    .X(\e1.alu1.out[26] ));
 sky130_fd_sc_hd__mux2_1 _13086_ (.A0(_00369_),
    .A1(\e1.alu1.a1.b[27] ),
    .S(net1),
    .X(\e1.alu1.out[27] ));
 sky130_fd_sc_hd__mux2_1 _13087_ (.A0(_00375_),
    .A1(\e1.alu1.a1.b[28] ),
    .S(net1),
    .X(\e1.alu1.out[28] ));
 sky130_fd_sc_hd__mux2_1 _13088_ (.A0(_00381_),
    .A1(\e1.alu1.a1.b[29] ),
    .S(net1),
    .X(\e1.alu1.out[29] ));
 sky130_fd_sc_hd__mux2_1 _13089_ (.A0(_00387_),
    .A1(\e1.alu1.a1.b[30] ),
    .S(net1),
    .X(\e1.alu1.out[30] ));
 sky130_fd_sc_hd__mux2_2 _13090_ (.A0(_00393_),
    .A1(\e1.alu1.a1.b[31] ),
    .S(net1),
    .X(\e1.alu1.out[31] ));
 sky130_fd_sc_hd__mux2_2 _13091_ (.A0(\next_pc[2] ),
    .A1(data_address[2]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _13092_ (.A0(\next_pc[3] ),
    .A1(data_address[3]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _13093_ (.A0(\next_pc[4] ),
    .A1(data_address[4]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _13094_ (.A0(\next_pc[5] ),
    .A1(data_address[5]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _13095_ (.A0(\next_pc[6] ),
    .A1(data_address[6]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _13096_ (.A0(\next_pc[7] ),
    .A1(data_address[7]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _13097_ (.A0(\next_pc[8] ),
    .A1(data_address[8]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _13098_ (.A0(\next_pc[9] ),
    .A1(data_address[9]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _13099_ (.A0(\next_pc[10] ),
    .A1(data_address[10]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _13100_ (.A0(\next_pc[11] ),
    .A1(data_address[11]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _13101_ (.A0(\next_pc[12] ),
    .A1(data_address[12]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _13102_ (.A0(\next_pc[13] ),
    .A1(data_address[13]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _13103_ (.A0(\next_pc[14] ),
    .A1(data_address[14]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _13104_ (.A0(\next_pc[15] ),
    .A1(data_address[15]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _13105_ (.A0(\next_pc[16] ),
    .A1(data_address[16]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _13106_ (.A0(\next_pc[17] ),
    .A1(data_address[17]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _13107_ (.A0(\next_pc[18] ),
    .A1(data_address[18]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _13108_ (.A0(\next_pc[19] ),
    .A1(data_address[19]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _13109_ (.A0(\next_pc[20] ),
    .A1(data_address[20]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _13110_ (.A0(\next_pc[21] ),
    .A1(data_address[21]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _13111_ (.A0(\next_pc[22] ),
    .A1(data_address[22]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _13112_ (.A0(\next_pc[23] ),
    .A1(data_address[23]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _13113_ (.A0(\next_pc[24] ),
    .A1(data_address[24]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _13114_ (.A0(\next_pc[25] ),
    .A1(data_address[25]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _13115_ (.A0(\next_pc[26] ),
    .A1(data_address[26]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _13116_ (.A0(\next_pc[27] ),
    .A1(data_address[27]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _13117_ (.A0(\next_pc[28] ),
    .A1(data_address[28]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _13118_ (.A0(\next_pc[29] ),
    .A1(data_address[29]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _13119_ (.A0(\next_pc[30] ),
    .A1(data_address[30]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _13120_ (.A0(\next_pc[31] ),
    .A1(data_address[31]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _13121_ (.A0(\e1.alu1.a[31] ),
    .A1(\e1.pc[31] ),
    .S(_00014_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_2 _13122_ (.A0(_00087_),
    .A1(_01270_),
    .S(_00014_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _13123_ (.A0(_00085_),
    .A1(_01268_),
    .S(_00014_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_2 _13124_ (.A0(_00084_),
    .A1(_01266_),
    .S(_00014_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _13125_ (.A0(_00081_),
    .A1(_01264_),
    .S(_00014_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _13126_ (.A0(_00080_),
    .A1(_01262_),
    .S(_00014_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _13127_ (.A0(_00078_),
    .A1(_01260_),
    .S(_00014_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _13128_ (.A0(_00077_),
    .A1(_01258_),
    .S(_00014_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _13129_ (.A0(_00073_),
    .A1(_01256_),
    .S(_00014_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _13130_ (.A0(_00072_),
    .A1(_01254_),
    .S(_00014_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _13131_ (.A0(_00070_),
    .A1(_01252_),
    .S(_00014_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_2 _13132_ (.A0(_00069_),
    .A1(_01250_),
    .S(_00014_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_2 _13133_ (.A0(_00066_),
    .A1(_01248_),
    .S(_00014_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _13134_ (.A0(_00065_),
    .A1(_01246_),
    .S(_00014_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _13135_ (.A0(_00063_),
    .A1(_01244_),
    .S(_00014_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _13136_ (.A0(_00062_),
    .A1(_01242_),
    .S(_00014_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _13137_ (.A0(_00057_),
    .A1(_01240_),
    .S(_00014_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _13138_ (.A0(_00056_),
    .A1(_01238_),
    .S(_00014_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _13139_ (.A0(_00054_),
    .A1(_01236_),
    .S(_00014_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _13140_ (.A0(_00053_),
    .A1(_01234_),
    .S(_00014_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_2 _13141_ (.A0(_00050_),
    .A1(_01232_),
    .S(_00014_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _13142_ (.A0(_00049_),
    .A1(_01230_),
    .S(_00014_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _13143_ (.A0(_00047_),
    .A1(_01228_),
    .S(_00014_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_2 _13144_ (.A0(_00046_),
    .A1(_01226_),
    .S(_00014_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _13145_ (.A0(_00042_),
    .A1(_01224_),
    .S(_00014_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_2 _13146_ (.A0(_00041_),
    .A1(_01222_),
    .S(_00014_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _13147_ (.A0(_00039_),
    .A1(_01220_),
    .S(_00014_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _13148_ (.A0(_00038_),
    .A1(_01218_),
    .S(_00014_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_2 _13149_ (.A0(_00035_),
    .A1(_01216_),
    .S(_00014_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_2 _13150_ (.A0(_00034_),
    .A1(_01214_),
    .S(_00014_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(_00032_),
    .A1(_01212_),
    .S(_00014_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _13152_ (.A0(_00031_),
    .A1(_01210_),
    .S(_00014_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _13153_ (.A0(_00407_),
    .A1(_00406_),
    .S(_00394_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _13154_ (.A0(_00404_),
    .A1(_00403_),
    .S(_00394_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _13155_ (.A0(_00401_),
    .A1(_00400_),
    .S(_00394_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _13156_ (.A0(_00398_),
    .A1(_00397_),
    .S(_00394_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _13157_ (.A0(_00395_),
    .A1(net50),
    .S(_00394_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _13158_ (.A0(_00088_),
    .A1(_00087_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _13159_ (.A0(_00388_),
    .A1(_00376_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _13160_ (.A0(_00389_),
    .A1(_00365_),
    .S(net9),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _13161_ (.A0(_00390_),
    .A1(_00342_),
    .S(net8),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_2 _13162_ (.A0(_00391_),
    .A1(_00296_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _13163_ (.A0(_00087_),
    .A1(_00085_),
    .S(net11),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _13164_ (.A0(_00382_),
    .A1(_00370_),
    .S(net10),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _13165_ (.A0(_00383_),
    .A1(_00359_),
    .S(net9),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _13166_ (.A0(_00384_),
    .A1(_00336_),
    .S(net8),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_2 _13167_ (.A0(_00385_),
    .A1(_00288_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _13168_ (.A0(_00376_),
    .A1(_00364_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _13169_ (.A0(_00377_),
    .A1(_00353_),
    .S(net9),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _13170_ (.A0(_00378_),
    .A1(_00330_),
    .S(net8),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _13171_ (.A0(_00379_),
    .A1(_00279_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _13172_ (.A0(_00085_),
    .A1(_00084_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _13173_ (.A0(_00370_),
    .A1(_00358_),
    .S(net10),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _13174_ (.A0(_00371_),
    .A1(_00347_),
    .S(net9),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _13175_ (.A0(_00372_),
    .A1(_00324_),
    .S(net8),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _13176_ (.A0(_00373_),
    .A1(_00270_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _13177_ (.A0(_00084_),
    .A1(_00081_),
    .S(net11),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _13178_ (.A0(_00365_),
    .A1(_00341_),
    .S(net9),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _13179_ (.A0(_00366_),
    .A1(_00318_),
    .S(net8),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _13180_ (.A0(_00367_),
    .A1(_00261_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _13181_ (.A0(_00364_),
    .A1(_00352_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _13182_ (.A0(_00081_),
    .A1(_00080_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _13183_ (.A0(_00359_),
    .A1(_00335_),
    .S(net9),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _13184_ (.A0(_00360_),
    .A1(_00312_),
    .S(net8),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _13185_ (.A0(_00361_),
    .A1(_00252_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _13186_ (.A0(_00358_),
    .A1(_00346_),
    .S(net10),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _13187_ (.A0(_00080_),
    .A1(_00078_),
    .S(net11),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _13188_ (.A0(_00353_),
    .A1(_00329_),
    .S(\e1.alu1.a1.b[2] ),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _13189_ (.A0(_00354_),
    .A1(_00306_),
    .S(net8),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _13190_ (.A0(_00355_),
    .A1(_00243_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _13191_ (.A0(_00352_),
    .A1(_00340_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _13192_ (.A0(_00078_),
    .A1(_00077_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _13193_ (.A0(_00347_),
    .A1(_00323_),
    .S(net9),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _13194_ (.A0(_00348_),
    .A1(_00300_),
    .S(net8),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _13195_ (.A0(_00349_),
    .A1(_00234_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _13196_ (.A0(_00346_),
    .A1(_00334_),
    .S(net10),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _13197_ (.A0(_00077_),
    .A1(_00073_),
    .S(net11),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _13198_ (.A0(_00342_),
    .A1(_00295_),
    .S(net8),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _13199_ (.A0(_00343_),
    .A1(_00225_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _13200_ (.A0(_00341_),
    .A1(_00317_),
    .S(net9),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _13201_ (.A0(_00340_),
    .A1(_00328_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _13202_ (.A0(_00073_),
    .A1(_00072_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _13203_ (.A0(_00336_),
    .A1(_00287_),
    .S(net8),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _13204_ (.A0(_00337_),
    .A1(_00213_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _13205_ (.A0(_00335_),
    .A1(_00311_),
    .S(net9),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _13206_ (.A0(_00334_),
    .A1(_00322_),
    .S(net10),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _13207_ (.A0(_00072_),
    .A1(_00070_),
    .S(net11),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _13208_ (.A0(_00330_),
    .A1(_00278_),
    .S(net8),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _13209_ (.A0(_00331_),
    .A1(_00200_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _13210_ (.A0(_00329_),
    .A1(_00305_),
    .S(\e1.alu1.a1.b[2] ),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _13211_ (.A0(_00328_),
    .A1(_00316_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _13212_ (.A0(_00070_),
    .A1(_00069_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _13213_ (.A0(_00324_),
    .A1(_00269_),
    .S(net8),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _13214_ (.A0(_00325_),
    .A1(_00187_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _13215_ (.A0(_00323_),
    .A1(_00299_),
    .S(net9),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _13216_ (.A0(_00322_),
    .A1(_00310_),
    .S(net10),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(_00069_),
    .A1(_00066_),
    .S(net11),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _13218_ (.A0(_00318_),
    .A1(_00260_),
    .S(net8),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(_00319_),
    .A1(_00174_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _13220_ (.A0(_00317_),
    .A1(_00294_),
    .S(net9),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(_00316_),
    .A1(_00304_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _13222_ (.A0(_00066_),
    .A1(_00065_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _13223_ (.A0(_00312_),
    .A1(_00251_),
    .S(net8),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _13224_ (.A0(_00313_),
    .A1(_00155_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _13225_ (.A0(_00311_),
    .A1(_00286_),
    .S(net9),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _13226_ (.A0(_00310_),
    .A1(_00298_),
    .S(net10),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _13227_ (.A0(_00065_),
    .A1(_00063_),
    .S(net11),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _13228_ (.A0(_00306_),
    .A1(_00242_),
    .S(\e1.alu1.a1.b[3] ),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _13229_ (.A0(_00307_),
    .A1(_00133_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _13230_ (.A0(_00305_),
    .A1(_00277_),
    .S(\e1.alu1.a1.b[2] ),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _13231_ (.A0(_00304_),
    .A1(_00293_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _13232_ (.A0(_00063_),
    .A1(_00062_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _13233_ (.A0(_00300_),
    .A1(_00233_),
    .S(net8),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_2 _13234_ (.A0(_00301_),
    .A1(_00095_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _13235_ (.A0(_00299_),
    .A1(_00268_),
    .S(net9),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _13236_ (.A0(_00298_),
    .A1(_00285_),
    .S(net10),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _13237_ (.A0(_00062_),
    .A1(_00057_),
    .S(net11),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_2 _13238_ (.A0(_00295_),
    .A1(_00224_),
    .S(net8),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _13239_ (.A0(_00294_),
    .A1(_00259_),
    .S(\e1.alu1.a1.b[2] ),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _13240_ (.A0(_00293_),
    .A1(_00276_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _13241_ (.A0(_00057_),
    .A1(_00056_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _13242_ (.A0(_00216_),
    .A1(_00218_),
    .S(net8),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _13243_ (.A0(_00290_),
    .A1(_00291_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_2 _13244_ (.A0(_00287_),
    .A1(_00284_),
    .S(net8),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _13245_ (.A0(_00286_),
    .A1(_00250_),
    .S(net9),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _13246_ (.A0(_00285_),
    .A1(_00267_),
    .S(net10),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _13247_ (.A0(_00056_),
    .A1(_00054_),
    .S(net11),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _13248_ (.A0(_00203_),
    .A1(_00205_),
    .S(net8),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _13249_ (.A0(_00281_),
    .A1(_00282_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_2 _13250_ (.A0(_00278_),
    .A1(_00275_),
    .S(net8),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _13251_ (.A0(_00277_),
    .A1(_00241_),
    .S(\e1.alu1.a1.b[2] ),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _13252_ (.A0(_00276_),
    .A1(_00258_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _13253_ (.A0(_00054_),
    .A1(_00053_),
    .S(net11),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _13254_ (.A0(_00190_),
    .A1(_00192_),
    .S(net8),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _13255_ (.A0(_00272_),
    .A1(_00273_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_2 _13256_ (.A0(_00269_),
    .A1(_00266_),
    .S(net8),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _13257_ (.A0(_00268_),
    .A1(_00232_),
    .S(net9),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _13258_ (.A0(_00267_),
    .A1(_00249_),
    .S(net10),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _13259_ (.A0(_00053_),
    .A1(_00050_),
    .S(net11),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _13260_ (.A0(_00177_),
    .A1(_00179_),
    .S(net8),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _13261_ (.A0(_00263_),
    .A1(_00264_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_2 _13262_ (.A0(_00260_),
    .A1(_00257_),
    .S(net8),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _13263_ (.A0(_00259_),
    .A1(_00223_),
    .S(\e1.alu1.a1.b[2] ),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _13264_ (.A0(_00258_),
    .A1(_00240_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _13265_ (.A0(_00050_),
    .A1(_00049_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _13266_ (.A0(_00162_),
    .A1(_00166_),
    .S(net8),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _13267_ (.A0(_00254_),
    .A1(_00255_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_2 _13268_ (.A0(_00251_),
    .A1(_00248_),
    .S(net8),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _13269_ (.A0(_00250_),
    .A1(_00210_),
    .S(net9),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _13270_ (.A0(_00249_),
    .A1(_00231_),
    .S(net10),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _13271_ (.A0(_00049_),
    .A1(_00047_),
    .S(net11),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _13272_ (.A0(_00142_),
    .A1(_00146_),
    .S(net8),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _13273_ (.A0(_00245_),
    .A1(_00246_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_2 _13274_ (.A0(_00242_),
    .A1(_00239_),
    .S(\e1.alu1.a1.b[3] ),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _13275_ (.A0(_00241_),
    .A1(_00197_),
    .S(\e1.alu1.a1.b[2] ),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _13276_ (.A0(_00240_),
    .A1(_00222_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _13277_ (.A0(_00047_),
    .A1(_00046_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _13278_ (.A0(_00113_),
    .A1(_00121_),
    .S(net8),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _13279_ (.A0(_00236_),
    .A1(_00237_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_2 _13280_ (.A0(_00233_),
    .A1(_00230_),
    .S(net8),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _13281_ (.A0(_00232_),
    .A1(_00184_),
    .S(net9),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _13282_ (.A0(_00231_),
    .A1(_00209_),
    .S(net10),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _13283_ (.A0(_00046_),
    .A1(_00042_),
    .S(net11),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _13284_ (.A0(_00060_),
    .A1(_00076_),
    .S(net8),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _13285_ (.A0(_00227_),
    .A1(_00228_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _13286_ (.A0(_00223_),
    .A1(_00173_),
    .S(\e1.alu1.a1.b[2] ),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _13287_ (.A0(_00222_),
    .A1(_00196_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _13288_ (.A0(_00042_),
    .A1(_00041_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _13289_ (.A0(_00158_),
    .A1(_00160_),
    .S(net9),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _13290_ (.A0(_00215_),
    .A1(_00216_),
    .S(net8),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _13291_ (.A0(_00217_),
    .A1(_00220_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _13292_ (.A0(_00218_),
    .A1(_00219_),
    .S(net8),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _13293_ (.A0(_00165_),
    .A1(_00167_),
    .S(net9),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _13294_ (.A0(_00161_),
    .A1(_00164_),
    .S(net9),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _13295_ (.A0(_00211_),
    .A1(_00154_),
    .S(net9),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _13296_ (.A0(_00209_),
    .A1(_00183_),
    .S(net10),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _13297_ (.A0(_00041_),
    .A1(_00039_),
    .S(net11),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _13298_ (.A0(_00138_),
    .A1(_00140_),
    .S(net9),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _13299_ (.A0(_00202_),
    .A1(_00203_),
    .S(net8),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _13300_ (.A0(_00204_),
    .A1(_00207_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_2 _13301_ (.A0(_00205_),
    .A1(_00206_),
    .S(net8),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _13302_ (.A0(_00145_),
    .A1(_00147_),
    .S(net9),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _13303_ (.A0(_00141_),
    .A1(_00144_),
    .S(net9),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _13304_ (.A0(_00198_),
    .A1(_00132_),
    .S(\e1.alu1.a1.b[2] ),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _13305_ (.A0(_00196_),
    .A1(_00172_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _13306_ (.A0(_00039_),
    .A1(_00038_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _13307_ (.A0(_00105_),
    .A1(_00109_),
    .S(net9),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _13308_ (.A0(_00189_),
    .A1(_00190_),
    .S(net8),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _13309_ (.A0(_00191_),
    .A1(_00194_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_2 _13310_ (.A0(_00192_),
    .A1(_00193_),
    .S(net8),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _13311_ (.A0(_00120_),
    .A1(_00124_),
    .S(net9),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _13312_ (.A0(_00112_),
    .A1(_00117_),
    .S(net9),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _13313_ (.A0(_00185_),
    .A1(_00094_),
    .S(net9),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _13314_ (.A0(_00183_),
    .A1(_00152_),
    .S(net10),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _13315_ (.A0(_00038_),
    .A1(_00035_),
    .S(net11),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _13316_ (.A0(_00044_),
    .A1(_00052_),
    .S(net9),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _13317_ (.A0(_00176_),
    .A1(_00177_),
    .S(net8),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _13318_ (.A0(_00178_),
    .A1(_00181_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _13319_ (.A0(_00179_),
    .A1(_00180_),
    .S(net8),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _13320_ (.A0(_00075_),
    .A1(_00083_),
    .S(net9),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _13321_ (.A0(_00059_),
    .A1(_00068_),
    .S(net9),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _13322_ (.A0(_00172_),
    .A1(_00131_),
    .S(\e1.alu1.a1.b[1] ),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _13323_ (.A0(_00035_),
    .A1(_00034_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _13324_ (.A0(_00101_),
    .A1(_00103_),
    .S(net10),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _13325_ (.A0(_00157_),
    .A1(_00158_),
    .S(net9),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _13326_ (.A0(_00159_),
    .A1(_00162_),
    .S(net8),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _13327_ (.A0(_00163_),
    .A1(_00170_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_2 _13328_ (.A0(_00166_),
    .A1(_00169_),
    .S(net8),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _13329_ (.A0(_00167_),
    .A1(_00168_),
    .S(net9),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _13330_ (.A0(_00123_),
    .A1(_00125_),
    .S(net10),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _13331_ (.A0(_00164_),
    .A1(_00165_),
    .S(net9),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _13332_ (.A0(_00119_),
    .A1(_00122_),
    .S(net10),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _13333_ (.A0(_00116_),
    .A1(_00118_),
    .S(net10),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _13334_ (.A0(_00160_),
    .A1(_00161_),
    .S(net9),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _13335_ (.A0(_00111_),
    .A1(_00115_),
    .S(net10),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _13336_ (.A0(_00108_),
    .A1(_00110_),
    .S(net10),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _13337_ (.A0(_00104_),
    .A1(_00107_),
    .S(net10),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _13338_ (.A0(_00153_),
    .A1(_00024_),
    .S(net10),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _13339_ (.A0(_00034_),
    .A1(_00032_),
    .S(net11),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _13340_ (.A0(_00036_),
    .A1(_00040_),
    .S(net10),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _13341_ (.A0(_00137_),
    .A1(_00138_),
    .S(net9),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _13342_ (.A0(_00139_),
    .A1(_00142_),
    .S(net8),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _13343_ (.A0(_00143_),
    .A1(_00150_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _13344_ (.A0(_00146_),
    .A1(_00149_),
    .S(net8),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _13345_ (.A0(_00147_),
    .A1(_00148_),
    .S(net9),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _13346_ (.A0(_00082_),
    .A1(_00086_),
    .S(net10),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _13347_ (.A0(_00144_),
    .A1(_00145_),
    .S(net9),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _13348_ (.A0(_00074_),
    .A1(_00079_),
    .S(net10),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _13349_ (.A0(_00067_),
    .A1(_00071_),
    .S(net10),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _13350_ (.A0(_00140_),
    .A1(_00141_),
    .S(net9),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _13351_ (.A0(_00058_),
    .A1(_00064_),
    .S(net10),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _13352_ (.A0(_00051_),
    .A1(_00055_),
    .S(net10),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _13353_ (.A0(_00043_),
    .A1(_00048_),
    .S(net10),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_2 _13354_ (.A0(_00134_),
    .A1(_00031_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _13355_ (.A0(_00032_),
    .A1(_00031_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _13356_ (.A0(_00032_),
    .A1(_00034_),
    .S(net11),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _13357_ (.A0(_00100_),
    .A1(_00101_),
    .S(net10),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _13358_ (.A0(_00102_),
    .A1(_00105_),
    .S(net9),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _13359_ (.A0(_00106_),
    .A1(_00113_),
    .S(net8),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _13360_ (.A0(_00114_),
    .A1(_00129_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_2 _13361_ (.A0(_00121_),
    .A1(_00128_),
    .S(net8),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _13362_ (.A0(_00124_),
    .A1(_00127_),
    .S(net9),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _13363_ (.A0(_00125_),
    .A1(_00126_),
    .S(net10),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _13364_ (.A0(_00085_),
    .A1(_00087_),
    .S(net11),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _13365_ (.A0(_00122_),
    .A1(_00123_),
    .S(net10),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _13366_ (.A0(_00081_),
    .A1(_00084_),
    .S(net11),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _13367_ (.A0(_00078_),
    .A1(_00080_),
    .S(net11),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _13368_ (.A0(_00117_),
    .A1(_00120_),
    .S(net9),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _13369_ (.A0(_00118_),
    .A1(_00119_),
    .S(net10),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _13370_ (.A0(_00073_),
    .A1(_00077_),
    .S(net11),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _13371_ (.A0(_00070_),
    .A1(_00072_),
    .S(net11),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _13372_ (.A0(_00115_),
    .A1(_00116_),
    .S(net10),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _13373_ (.A0(_00066_),
    .A1(_00069_),
    .S(net11),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _13374_ (.A0(_00063_),
    .A1(_00065_),
    .S(net11),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _13375_ (.A0(_00109_),
    .A1(_00112_),
    .S(net9),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _13376_ (.A0(_00110_),
    .A1(_00111_),
    .S(net10),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _13377_ (.A0(_00057_),
    .A1(_00062_),
    .S(net11),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _13378_ (.A0(_00054_),
    .A1(_00056_),
    .S(net11),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _13379_ (.A0(_00107_),
    .A1(_00108_),
    .S(net10),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _13380_ (.A0(_00050_),
    .A1(_00053_),
    .S(net11),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _13381_ (.A0(_00047_),
    .A1(_00049_),
    .S(net11),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _13382_ (.A0(_00103_),
    .A1(_00104_),
    .S(net10),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _13383_ (.A0(_00042_),
    .A1(_00046_),
    .S(net11),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _13384_ (.A0(_00039_),
    .A1(_00041_),
    .S(net11),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _13385_ (.A0(_00035_),
    .A1(_00038_),
    .S(net11),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _13386_ (.A0(_00010_),
    .A1(_00005_),
    .S(_00097_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _13387_ (.A0(_00004_),
    .A1(\c1.instruction2[13] ),
    .S(\c1.instruction2[12] ),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _13388_ (.A0(_00031_),
    .A1(_00032_),
    .S(net11),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _13389_ (.A0(_00033_),
    .A1(_00036_),
    .S(net10),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _13390_ (.A0(_00037_),
    .A1(_00044_),
    .S(net9),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _13391_ (.A0(_00045_),
    .A1(_00060_),
    .S(net8),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_2 _13392_ (.A0(_00061_),
    .A1(_00092_),
    .S(\e1.alu1.a1.b[4] ),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _13393_ (.A0(_00076_),
    .A1(_00091_),
    .S(net8),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _13394_ (.A0(_00083_),
    .A1(_00090_),
    .S(net9),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _13395_ (.A0(_00086_),
    .A1(_00089_),
    .S(net10),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _13396_ (.A0(_00087_),
    .A1(_00088_),
    .S(\e1.alu1.a1.b[0] ),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _13397_ (.A0(_00084_),
    .A1(_00085_),
    .S(net11),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _13398_ (.A0(_00079_),
    .A1(_00082_),
    .S(net10),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _13399_ (.A0(_00080_),
    .A1(_00081_),
    .S(net11),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _13400_ (.A0(_00077_),
    .A1(_00078_),
    .S(net11),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _13401_ (.A0(_00068_),
    .A1(_00075_),
    .S(net9),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _13402_ (.A0(_00071_),
    .A1(_00074_),
    .S(net10),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _13403_ (.A0(_00072_),
    .A1(_00073_),
    .S(net11),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _13404_ (.A0(_00069_),
    .A1(_00070_),
    .S(net11),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _13405_ (.A0(_00064_),
    .A1(_00067_),
    .S(net10),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _13406_ (.A0(_00065_),
    .A1(_00066_),
    .S(net11),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _13407_ (.A0(_00062_),
    .A1(_00063_),
    .S(net11),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _13408_ (.A0(_00052_),
    .A1(_00059_),
    .S(net9),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _13409_ (.A0(_00055_),
    .A1(_00058_),
    .S(net10),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _13410_ (.A0(_00056_),
    .A1(_00057_),
    .S(net11),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _13411_ (.A0(_00053_),
    .A1(_00054_),
    .S(net11),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _13412_ (.A0(_00048_),
    .A1(_00051_),
    .S(net10),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _13413_ (.A0(_00049_),
    .A1(_00050_),
    .S(net11),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _13414_ (.A0(_00046_),
    .A1(_00047_),
    .S(net11),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _13415_ (.A0(_00040_),
    .A1(_00043_),
    .S(net10),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _13416_ (.A0(_00041_),
    .A1(_00042_),
    .S(net11),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _13417_ (.A0(_00038_),
    .A1(_00039_),
    .S(net11),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _13418_ (.A0(_00034_),
    .A1(_00035_),
    .S(net11),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _13419_ (.A0(_00029_),
    .A1(_00021_),
    .S(_00022_),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _13420_ (.A0(_00009_),
    .A1(_00016_),
    .S(_00027_),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _13421_ (.A0(_00023_),
    .A1(_00008_),
    .S(_00025_),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _13422_ (.A0(_00006_),
    .A1(_00010_),
    .S(_00007_),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _13423_ (.A0(_00017_),
    .A1(_00012_),
    .S(_00007_),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _13424_ (.A0(\c1.instruction2[13] ),
    .A1(\c1.instruction2[14] ),
    .S(\c1.instruction2[12] ),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _13425_ (.A0(_00011_),
    .A1(_00012_),
    .S(_00007_),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _13426_ (.A0(\next_pc[1] ),
    .A1(data_address[1]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _13427_ (.A0(\next_pc[0] ),
    .A1(data_address[0]),
    .S(MEM_X_BRANCH_TAKEN),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _13428_ (.A0(_01202_),
    .A1(_01207_),
    .S(net54),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _13429_ (.A0(_01208_),
    .A1(rdata[31]),
    .S(\DEP_PLACE[2] ),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _13430_ (.A0(_01209_),
    .A1(\e1.alu1.out[31] ),
    .S(\DEP_PLACE[0] ),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _13431_ (.A0(_01190_),
    .A1(_01195_),
    .S(net54),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _13432_ (.A0(_01196_),
    .A1(rdata[30]),
    .S(net2),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _13433_ (.A0(_01197_),
    .A1(\e1.alu1.out[30] ),
    .S(\DEP_PLACE[0] ),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _13434_ (.A0(_01178_),
    .A1(_01183_),
    .S(net54),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _13435_ (.A0(_01184_),
    .A1(rdata[29]),
    .S(net2),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _13436_ (.A0(_01185_),
    .A1(\e1.alu1.out[29] ),
    .S(\DEP_PLACE[0] ),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _13437_ (.A0(_01166_),
    .A1(_01171_),
    .S(\c1.instruction1[19] ),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _13438_ (.A0(_01172_),
    .A1(rdata[28]),
    .S(net2),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _13439_ (.A0(_01173_),
    .A1(\e1.alu1.out[28] ),
    .S(\DEP_PLACE[0] ),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _13440_ (.A0(_01154_),
    .A1(_01159_),
    .S(\c1.instruction1[19] ),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _13441_ (.A0(_01160_),
    .A1(rdata[27]),
    .S(net2),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _13442_ (.A0(_01161_),
    .A1(\e1.alu1.out[27] ),
    .S(\DEP_PLACE[0] ),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _13443_ (.A0(_01142_),
    .A1(_01147_),
    .S(\c1.instruction1[19] ),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _13444_ (.A0(_01148_),
    .A1(rdata[26]),
    .S(net2),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _13445_ (.A0(_01149_),
    .A1(\e1.alu1.out[26] ),
    .S(\DEP_PLACE[0] ),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_2 _13446_ (.A0(_01130_),
    .A1(_01135_),
    .S(\c1.instruction1[19] ),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _13447_ (.A0(_01136_),
    .A1(rdata[25]),
    .S(net2),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _13448_ (.A0(_01137_),
    .A1(\e1.alu1.out[25] ),
    .S(\DEP_PLACE[0] ),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _13449_ (.A0(_01118_),
    .A1(_01123_),
    .S(\c1.instruction1[19] ),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_2 _13450_ (.A0(_01124_),
    .A1(rdata[24]),
    .S(net2),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _13451_ (.A0(_01125_),
    .A1(\e1.alu1.out[24] ),
    .S(\DEP_PLACE[0] ),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_2 _13452_ (.A0(_01106_),
    .A1(_01111_),
    .S(\c1.instruction1[19] ),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _13453_ (.A0(_01112_),
    .A1(rdata[23]),
    .S(net2),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _13454_ (.A0(_01113_),
    .A1(\e1.alu1.out[23] ),
    .S(\DEP_PLACE[0] ),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _13455_ (.A0(_01094_),
    .A1(_01099_),
    .S(net54),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_2 _13456_ (.A0(_01100_),
    .A1(rdata[22]),
    .S(net2),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _13457_ (.A0(_01101_),
    .A1(\e1.alu1.out[22] ),
    .S(\DEP_PLACE[0] ),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _13458_ (.A0(_01082_),
    .A1(_01087_),
    .S(net54),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_2 _13459_ (.A0(_01088_),
    .A1(rdata[21]),
    .S(net2),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _13460_ (.A0(_01089_),
    .A1(\e1.alu1.out[21] ),
    .S(\DEP_PLACE[0] ),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _13461_ (.A0(_01070_),
    .A1(_01075_),
    .S(net54),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_4 _13462_ (.A0(_01076_),
    .A1(rdata[20]),
    .S(net2),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _13463_ (.A0(_01077_),
    .A1(\e1.alu1.out[20] ),
    .S(\DEP_PLACE[0] ),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _13464_ (.A0(_01058_),
    .A1(_01063_),
    .S(net54),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_2 _13465_ (.A0(_01064_),
    .A1(rdata[19]),
    .S(net2),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _13466_ (.A0(_01065_),
    .A1(\e1.alu1.out[19] ),
    .S(\DEP_PLACE[0] ),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _13467_ (.A0(_01046_),
    .A1(_01051_),
    .S(net54),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _13468_ (.A0(_01052_),
    .A1(rdata[18]),
    .S(\DEP_PLACE[2] ),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _13469_ (.A0(_01053_),
    .A1(\e1.alu1.out[18] ),
    .S(\DEP_PLACE[0] ),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _13470_ (.A0(_01034_),
    .A1(_01039_),
    .S(net54),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _13471_ (.A0(_01040_),
    .A1(rdata[17]),
    .S(net2),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _13472_ (.A0(_01041_),
    .A1(\e1.alu1.out[17] ),
    .S(\DEP_PLACE[0] ),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _13473_ (.A0(_01022_),
    .A1(_01027_),
    .S(net54),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_2 _13474_ (.A0(_01028_),
    .A1(rdata[16]),
    .S(net2),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _13475_ (.A0(_01029_),
    .A1(\e1.alu1.out[16] ),
    .S(\DEP_PLACE[0] ),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_2 _13476_ (.A0(_01010_),
    .A1(_01015_),
    .S(net54),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _13477_ (.A0(_01016_),
    .A1(rdata[15]),
    .S(net2),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _13478_ (.A0(_01017_),
    .A1(\e1.alu1.out[15] ),
    .S(\DEP_PLACE[0] ),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _13479_ (.A0(_00998_),
    .A1(_01003_),
    .S(net54),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _13480_ (.A0(_01004_),
    .A1(rdata[14]),
    .S(net2),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _13481_ (.A0(_01005_),
    .A1(\e1.alu1.out[14] ),
    .S(\DEP_PLACE[0] ),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_2 _13482_ (.A0(_00986_),
    .A1(_00991_),
    .S(net54),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_2 _13483_ (.A0(_00992_),
    .A1(rdata[13]),
    .S(net2),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _13484_ (.A0(_00993_),
    .A1(\e1.alu1.out[13] ),
    .S(\DEP_PLACE[0] ),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_2 _13485_ (.A0(_00974_),
    .A1(_00979_),
    .S(net54),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _13486_ (.A0(_00980_),
    .A1(rdata[12]),
    .S(net2),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _13487_ (.A0(_00981_),
    .A1(\e1.alu1.out[12] ),
    .S(\DEP_PLACE[0] ),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _13488_ (.A0(_00962_),
    .A1(_00967_),
    .S(net54),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_2 _13489_ (.A0(_00968_),
    .A1(rdata[11]),
    .S(net2),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _13490_ (.A0(_00969_),
    .A1(\e1.alu1.out[11] ),
    .S(\DEP_PLACE[0] ),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_4 _13491_ (.A0(_00950_),
    .A1(_00955_),
    .S(net54),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _13492_ (.A0(_00956_),
    .A1(rdata[10]),
    .S(net2),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _13493_ (.A0(_00957_),
    .A1(\e1.alu1.out[10] ),
    .S(\DEP_PLACE[0] ),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_2 _13494_ (.A0(_00938_),
    .A1(_00943_),
    .S(net54),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_2 _13495_ (.A0(_00944_),
    .A1(rdata[9]),
    .S(net2),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _13496_ (.A0(_00945_),
    .A1(\e1.alu1.out[9] ),
    .S(\DEP_PLACE[0] ),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _13497_ (.A0(_00926_),
    .A1(_00931_),
    .S(net54),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_4 _13498_ (.A0(_00932_),
    .A1(rdata[8]),
    .S(net2),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _13499_ (.A0(_00933_),
    .A1(\e1.alu1.out[8] ),
    .S(\DEP_PLACE[0] ),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _13500_ (.A0(_00914_),
    .A1(_00919_),
    .S(net54),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_2 _13501_ (.A0(_00920_),
    .A1(rdata[7]),
    .S(net2),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _13502_ (.A0(_00921_),
    .A1(\e1.alu1.out[7] ),
    .S(\DEP_PLACE[0] ),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _13503_ (.A0(_00902_),
    .A1(_00907_),
    .S(net54),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_2 _13504_ (.A0(_00908_),
    .A1(rdata[6]),
    .S(net2),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _13505_ (.A0(_00909_),
    .A1(\e1.alu1.out[6] ),
    .S(\DEP_PLACE[0] ),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_4 _13506_ (.A0(_00890_),
    .A1(_00895_),
    .S(net54),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _13507_ (.A0(_00896_),
    .A1(rdata[5]),
    .S(\DEP_PLACE[2] ),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _13508_ (.A0(_00897_),
    .A1(\e1.alu1.out[5] ),
    .S(\DEP_PLACE[0] ),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_2 _13509_ (.A0(_00878_),
    .A1(_00883_),
    .S(net54),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _13510_ (.A0(_00884_),
    .A1(rdata[4]),
    .S(\DEP_PLACE[2] ),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _13511_ (.A0(_00885_),
    .A1(\e1.alu1.out[4] ),
    .S(\DEP_PLACE[0] ),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_2 _13512_ (.A0(_00866_),
    .A1(_00871_),
    .S(net54),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _13513_ (.A0(_00872_),
    .A1(rdata[3]),
    .S(\DEP_PLACE[2] ),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _13514_ (.A0(_00873_),
    .A1(\e1.alu1.out[3] ),
    .S(\DEP_PLACE[0] ),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _13515_ (.A0(_00854_),
    .A1(_00859_),
    .S(net54),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_2 _13516_ (.A0(_00860_),
    .A1(rdata[2]),
    .S(net2),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _13517_ (.A0(_00861_),
    .A1(\e1.alu1.out[2] ),
    .S(\DEP_PLACE[0] ),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _13518_ (.A0(_00842_),
    .A1(_00847_),
    .S(net54),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _13519_ (.A0(_00848_),
    .A1(rdata[1]),
    .S(\DEP_PLACE[2] ),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _13520_ (.A0(_00849_),
    .A1(\e1.alu1.out[1] ),
    .S(\DEP_PLACE[0] ),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _13521_ (.A0(_00830_),
    .A1(_00835_),
    .S(net54),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _13522_ (.A0(_00836_),
    .A1(rdata[0]),
    .S(\DEP_PLACE[2] ),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _13523_ (.A0(_00837_),
    .A1(\e1.alu1.out[0] ),
    .S(\DEP_PLACE[0] ),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _13524_ (.A0(_00817_),
    .A1(_00822_),
    .S(net53),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _13525_ (.A0(_00823_),
    .A1(net3),
    .S(_00420_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _13526_ (.A0(_00824_),
    .A1(\wbmemout[31] ),
    .S(\DEP_PLACE[3] ),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _13527_ (.A0(_00825_),
    .A1(\e1.alu1.out[31] ),
    .S(\DEP_PLACE[1] ),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _13528_ (.A0(_00804_),
    .A1(_00809_),
    .S(net53),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _13529_ (.A0(_00810_),
    .A1(net3),
    .S(net4),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _13530_ (.A0(_00811_),
    .A1(\wbmemout[30] ),
    .S(\DEP_PLACE[3] ),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _13531_ (.A0(_00812_),
    .A1(\e1.alu1.out[30] ),
    .S(\DEP_PLACE[1] ),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _13532_ (.A0(_00791_),
    .A1(_00796_),
    .S(net53),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _13533_ (.A0(_00797_),
    .A1(net3),
    .S(net4),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _13534_ (.A0(_00798_),
    .A1(\wbmemout[29] ),
    .S(\DEP_PLACE[3] ),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _13535_ (.A0(_00799_),
    .A1(\e1.alu1.out[29] ),
    .S(\DEP_PLACE[1] ),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _13536_ (.A0(_00778_),
    .A1(_00783_),
    .S(\c1.instruction1[24] ),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _13537_ (.A0(_00784_),
    .A1(net3),
    .S(net4),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _13538_ (.A0(_00785_),
    .A1(\wbmemout[28] ),
    .S(\DEP_PLACE[3] ),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _13539_ (.A0(_00786_),
    .A1(\e1.alu1.out[28] ),
    .S(\DEP_PLACE[1] ),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _13540_ (.A0(_00765_),
    .A1(_00770_),
    .S(\c1.instruction1[24] ),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _13541_ (.A0(_00771_),
    .A1(net3),
    .S(net4),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _13542_ (.A0(_00772_),
    .A1(\wbmemout[27] ),
    .S(\DEP_PLACE[3] ),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _13543_ (.A0(_00773_),
    .A1(\e1.alu1.out[27] ),
    .S(\DEP_PLACE[1] ),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _13544_ (.A0(_00752_),
    .A1(_00757_),
    .S(\c1.instruction1[24] ),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _13545_ (.A0(_00758_),
    .A1(net3),
    .S(net4),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _13546_ (.A0(_00759_),
    .A1(\wbmemout[26] ),
    .S(\DEP_PLACE[3] ),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _13547_ (.A0(_00760_),
    .A1(\e1.alu1.out[26] ),
    .S(\DEP_PLACE[1] ),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _13548_ (.A0(_00739_),
    .A1(_00744_),
    .S(\c1.instruction1[24] ),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _13549_ (.A0(_00745_),
    .A1(net3),
    .S(net4),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _13550_ (.A0(_00746_),
    .A1(\wbmemout[25] ),
    .S(\DEP_PLACE[3] ),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _13551_ (.A0(_00747_),
    .A1(\e1.alu1.out[25] ),
    .S(\DEP_PLACE[1] ),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _13552_ (.A0(_00726_),
    .A1(_00731_),
    .S(\c1.instruction1[24] ),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _13553_ (.A0(_00732_),
    .A1(net3),
    .S(net4),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_2 _13554_ (.A0(_00733_),
    .A1(\wbmemout[24] ),
    .S(\DEP_PLACE[3] ),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _13555_ (.A0(_00734_),
    .A1(\e1.alu1.out[24] ),
    .S(\DEP_PLACE[1] ),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_2 _13556_ (.A0(_00713_),
    .A1(_00718_),
    .S(\c1.instruction1[24] ),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _13557_ (.A0(_00719_),
    .A1(net3),
    .S(net4),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _13558_ (.A0(_00720_),
    .A1(\wbmemout[23] ),
    .S(\DEP_PLACE[3] ),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _13559_ (.A0(_00721_),
    .A1(\e1.alu1.out[23] ),
    .S(\DEP_PLACE[1] ),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _13560_ (.A0(_00700_),
    .A1(_00705_),
    .S(net53),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _13561_ (.A0(_00706_),
    .A1(net3),
    .S(net4),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_2 _13562_ (.A0(_00707_),
    .A1(\wbmemout[22] ),
    .S(\DEP_PLACE[3] ),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _13563_ (.A0(_00708_),
    .A1(\e1.alu1.out[22] ),
    .S(\DEP_PLACE[1] ),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _13564_ (.A0(_00687_),
    .A1(_00692_),
    .S(net53),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _13565_ (.A0(_00693_),
    .A1(net3),
    .S(net4),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_2 _13566_ (.A0(_00694_),
    .A1(\wbmemout[21] ),
    .S(\DEP_PLACE[3] ),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _13567_ (.A0(_00695_),
    .A1(\e1.alu1.out[21] ),
    .S(\DEP_PLACE[1] ),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _13568_ (.A0(_00674_),
    .A1(_00679_),
    .S(net53),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _13569_ (.A0(_00680_),
    .A1(net3),
    .S(net4),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_2 _13570_ (.A0(_00681_),
    .A1(\wbmemout[20] ),
    .S(\DEP_PLACE[3] ),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _13571_ (.A0(_00682_),
    .A1(\e1.alu1.out[20] ),
    .S(\DEP_PLACE[1] ),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _13572_ (.A0(_00661_),
    .A1(_00666_),
    .S(net53),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _13573_ (.A0(_00667_),
    .A1(net3),
    .S(net5),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_2 _13574_ (.A0(_00668_),
    .A1(\wbmemout[19] ),
    .S(\DEP_PLACE[3] ),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _13575_ (.A0(_00669_),
    .A1(\e1.alu1.out[19] ),
    .S(\DEP_PLACE[1] ),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _13576_ (.A0(_00648_),
    .A1(_00653_),
    .S(net53),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _13577_ (.A0(_00654_),
    .A1(net3),
    .S(_00420_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _13578_ (.A0(_00655_),
    .A1(\wbmemout[18] ),
    .S(\DEP_PLACE[3] ),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _13579_ (.A0(_00656_),
    .A1(\e1.alu1.out[18] ),
    .S(\DEP_PLACE[1] ),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _13580_ (.A0(_00635_),
    .A1(_00640_),
    .S(net53),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _13581_ (.A0(_00641_),
    .A1(net3),
    .S(net5),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _13582_ (.A0(_00642_),
    .A1(\wbmemout[17] ),
    .S(\DEP_PLACE[3] ),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _13583_ (.A0(_00643_),
    .A1(\e1.alu1.out[17] ),
    .S(\DEP_PLACE[1] ),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _13584_ (.A0(_00622_),
    .A1(_00627_),
    .S(net53),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _13585_ (.A0(_00628_),
    .A1(\d1.addr[11] ),
    .S(_00420_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _13586_ (.A0(_00629_),
    .A1(\wbmemout[16] ),
    .S(\DEP_PLACE[3] ),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _13587_ (.A0(_00630_),
    .A1(\e1.alu1.out[16] ),
    .S(\DEP_PLACE[1] ),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _13588_ (.A0(_00609_),
    .A1(_00614_),
    .S(net53),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _13589_ (.A0(_00615_),
    .A1(\d1.addr[11] ),
    .S(_00420_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _13590_ (.A0(_00616_),
    .A1(\wbmemout[15] ),
    .S(\DEP_PLACE[3] ),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _13591_ (.A0(_00617_),
    .A1(\e1.alu1.out[15] ),
    .S(\DEP_PLACE[1] ),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _13592_ (.A0(_00596_),
    .A1(_00601_),
    .S(net53),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _13593_ (.A0(_00602_),
    .A1(\d1.addr[11] ),
    .S(_00420_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _13594_ (.A0(_00603_),
    .A1(\wbmemout[14] ),
    .S(\DEP_PLACE[3] ),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _13595_ (.A0(_00604_),
    .A1(\e1.alu1.out[14] ),
    .S(\DEP_PLACE[1] ),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_2 _13596_ (.A0(_00583_),
    .A1(_00588_),
    .S(net53),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _13597_ (.A0(_00589_),
    .A1(\d1.addr[11] ),
    .S(_00420_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _13598_ (.A0(_00590_),
    .A1(\wbmemout[13] ),
    .S(\DEP_PLACE[3] ),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _13599_ (.A0(_00591_),
    .A1(\e1.alu1.out[13] ),
    .S(\DEP_PLACE[1] ),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_2 _13600_ (.A0(_00570_),
    .A1(_00575_),
    .S(net53),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _13601_ (.A0(_00576_),
    .A1(\d1.addr[11] ),
    .S(_00420_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _13602_ (.A0(_00577_),
    .A1(\wbmemout[12] ),
    .S(\DEP_PLACE[3] ),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _13603_ (.A0(_00578_),
    .A1(\e1.alu1.out[12] ),
    .S(\DEP_PLACE[1] ),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_2 _13604_ (.A0(_00557_),
    .A1(_00562_),
    .S(net53),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _13605_ (.A0(_00563_),
    .A1(\d1.addr[11] ),
    .S(_00420_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _13606_ (.A0(_00564_),
    .A1(\wbmemout[11] ),
    .S(\DEP_PLACE[3] ),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _13607_ (.A0(_00565_),
    .A1(\e1.alu1.out[11] ),
    .S(\DEP_PLACE[1] ),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_4 _13608_ (.A0(_00544_),
    .A1(_00549_),
    .S(net53),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _13609_ (.A0(_00550_),
    .A1(\d1.addr[10] ),
    .S(_00420_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _13610_ (.A0(_00551_),
    .A1(\wbmemout[10] ),
    .S(\DEP_PLACE[3] ),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _13611_ (.A0(_00552_),
    .A1(\e1.alu1.out[10] ),
    .S(\DEP_PLACE[1] ),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_4 _13612_ (.A0(_00531_),
    .A1(_00536_),
    .S(net53),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _13613_ (.A0(_00537_),
    .A1(\d1.addr[9] ),
    .S(_00420_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _13614_ (.A0(_00538_),
    .A1(\wbmemout[9] ),
    .S(\DEP_PLACE[3] ),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _13615_ (.A0(_00539_),
    .A1(\e1.alu1.out[9] ),
    .S(\DEP_PLACE[1] ),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_2 _13616_ (.A0(_00518_),
    .A1(_00523_),
    .S(net53),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _13617_ (.A0(_00524_),
    .A1(\d1.addr[8] ),
    .S(net5),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _13618_ (.A0(_00525_),
    .A1(\wbmemout[8] ),
    .S(\DEP_PLACE[3] ),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _13619_ (.A0(_00526_),
    .A1(\e1.alu1.out[8] ),
    .S(\DEP_PLACE[1] ),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_2 _13620_ (.A0(_00505_),
    .A1(_00510_),
    .S(net53),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _13621_ (.A0(_00511_),
    .A1(\d1.addr[7] ),
    .S(net5),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_2 _13622_ (.A0(_00512_),
    .A1(\wbmemout[7] ),
    .S(\DEP_PLACE[3] ),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _13623_ (.A0(_00513_),
    .A1(\e1.alu1.out[7] ),
    .S(\DEP_PLACE[1] ),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_2 _13624_ (.A0(_00492_),
    .A1(_00497_),
    .S(net53),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _13625_ (.A0(_00498_),
    .A1(\d1.addr[6] ),
    .S(net5),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_2 _13626_ (.A0(_00499_),
    .A1(\wbmemout[6] ),
    .S(\DEP_PLACE[3] ),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _13627_ (.A0(_00500_),
    .A1(\e1.alu1.out[6] ),
    .S(\DEP_PLACE[1] ),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_2 _13628_ (.A0(_00479_),
    .A1(_00484_),
    .S(net53),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _13629_ (.A0(_00485_),
    .A1(\d1.addr[5] ),
    .S(net5),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _13630_ (.A0(_00486_),
    .A1(\wbmemout[5] ),
    .S(\DEP_PLACE[3] ),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _13631_ (.A0(_00487_),
    .A1(\e1.alu1.out[5] ),
    .S(\DEP_PLACE[1] ),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_2 _13632_ (.A0(_00466_),
    .A1(_00471_),
    .S(net53),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _13633_ (.A0(_00472_),
    .A1(\d1.addr[4] ),
    .S(net5),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _13634_ (.A0(_00473_),
    .A1(\wbmemout[4] ),
    .S(\DEP_PLACE[3] ),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _13635_ (.A0(_00474_),
    .A1(\e1.alu1.out[4] ),
    .S(\DEP_PLACE[1] ),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_2 _13636_ (.A0(_00453_),
    .A1(_00458_),
    .S(net53),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _13637_ (.A0(_00459_),
    .A1(\d1.addr[3] ),
    .S(net5),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _13638_ (.A0(_00460_),
    .A1(\wbmemout[3] ),
    .S(\DEP_PLACE[3] ),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _13639_ (.A0(_00461_),
    .A1(\e1.alu1.out[3] ),
    .S(\DEP_PLACE[1] ),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_2 _13640_ (.A0(_00440_),
    .A1(_00445_),
    .S(net53),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _13641_ (.A0(_00446_),
    .A1(\d1.addr[2] ),
    .S(net5),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _13642_ (.A0(_00447_),
    .A1(\wbmemout[2] ),
    .S(\DEP_PLACE[3] ),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _13643_ (.A0(_00448_),
    .A1(\e1.alu1.out[2] ),
    .S(\DEP_PLACE[1] ),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _13644_ (.A0(_00427_),
    .A1(_00432_),
    .S(net53),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _13645_ (.A0(_00433_),
    .A1(\d1.addr[1] ),
    .S(_00420_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _13646_ (.A0(_00434_),
    .A1(\wbmemout[1] ),
    .S(\DEP_PLACE[3] ),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _13647_ (.A0(_00435_),
    .A1(\e1.alu1.out[1] ),
    .S(\DEP_PLACE[1] ),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _13648_ (.A0(_00413_),
    .A1(_00418_),
    .S(net53),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _13649_ (.A0(_00419_),
    .A1(\d1.addr[0] ),
    .S(_00420_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _13650_ (.A0(_00421_),
    .A1(\wbmemout[0] ),
    .S(\DEP_PLACE[3] ),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _13651_ (.A0(_00422_),
    .A1(\e1.alu1.out[0] ),
    .S(\DEP_PLACE[1] ),
    .X(_01273_));
 sky130_fd_sc_hd__mux4_1 _13652_ (.A0(\r1.regblock[0][31] ),
    .A1(\r1.regblock[1][31] ),
    .A2(\r1.regblock[2][31] ),
    .A3(\r1.regblock[3][31] ),
    .S0(net27),
    .S1(net20),
    .X(_01198_));
 sky130_fd_sc_hd__mux4_2 _13653_ (.A0(\r1.regblock[4][31] ),
    .A1(\r1.regblock[5][31] ),
    .A2(\r1.regblock[6][31] ),
    .A3(\r1.regblock[7][31] ),
    .S0(net25),
    .S1(net18),
    .X(_01199_));
 sky130_fd_sc_hd__mux4_1 _13654_ (.A0(\r1.regblock[8][31] ),
    .A1(\r1.regblock[9][31] ),
    .A2(\r1.regblock[10][31] ),
    .A3(\r1.regblock[11][31] ),
    .S0(net27),
    .S1(net20),
    .X(_01200_));
 sky130_fd_sc_hd__mux4_1 _13655_ (.A0(\r1.regblock[12][31] ),
    .A1(\r1.regblock[13][31] ),
    .A2(\r1.regblock[14][31] ),
    .A3(\r1.regblock[15][31] ),
    .S0(net27),
    .S1(net20),
    .X(_01201_));
 sky130_fd_sc_hd__mux4_2 _13656_ (.A0(_01198_),
    .A1(_01199_),
    .A2(_01200_),
    .A3(_01201_),
    .S0(net14),
    .S1(net12),
    .X(_01202_));
 sky130_fd_sc_hd__mux4_2 _13657_ (.A0(\r1.regblock[16][31] ),
    .A1(\r1.regblock[17][31] ),
    .A2(\r1.regblock[18][31] ),
    .A3(\r1.regblock[19][31] ),
    .S0(net28),
    .S1(net20),
    .X(_01203_));
 sky130_fd_sc_hd__mux4_1 _13658_ (.A0(\r1.regblock[20][31] ),
    .A1(\r1.regblock[21][31] ),
    .A2(\r1.regblock[22][31] ),
    .A3(\r1.regblock[23][31] ),
    .S0(net28),
    .S1(net20),
    .X(_01204_));
 sky130_fd_sc_hd__mux4_1 _13659_ (.A0(\r1.regblock[24][31] ),
    .A1(\r1.regblock[25][31] ),
    .A2(\r1.regblock[26][31] ),
    .A3(\r1.regblock[27][31] ),
    .S0(net28),
    .S1(net20),
    .X(_01205_));
 sky130_fd_sc_hd__mux4_2 _13660_ (.A0(\r1.regblock[28][31] ),
    .A1(\r1.regblock[29][31] ),
    .A2(\r1.regblock[30][31] ),
    .A3(\r1.regblock[31][31] ),
    .S0(net27),
    .S1(net20),
    .X(_01206_));
 sky130_fd_sc_hd__mux4_1 _13661_ (.A0(_01203_),
    .A1(_01204_),
    .A2(_01205_),
    .A3(_01206_),
    .S0(net15),
    .S1(\c1.instruction1[18] ),
    .X(_01207_));
 sky130_fd_sc_hd__mux4_1 _13662_ (.A0(\r1.regblock[0][30] ),
    .A1(\r1.regblock[1][30] ),
    .A2(\r1.regblock[2][30] ),
    .A3(\r1.regblock[3][30] ),
    .S0(net27),
    .S1(net20),
    .X(_01186_));
 sky130_fd_sc_hd__mux4_2 _13663_ (.A0(\r1.regblock[4][30] ),
    .A1(\r1.regblock[5][30] ),
    .A2(\r1.regblock[6][30] ),
    .A3(\r1.regblock[7][30] ),
    .S0(net27),
    .S1(net19),
    .X(_01187_));
 sky130_fd_sc_hd__mux4_2 _13664_ (.A0(\r1.regblock[8][30] ),
    .A1(\r1.regblock[9][30] ),
    .A2(\r1.regblock[10][30] ),
    .A3(\r1.regblock[11][30] ),
    .S0(net27),
    .S1(net20),
    .X(_01188_));
 sky130_fd_sc_hd__mux4_1 _13665_ (.A0(\r1.regblock[12][30] ),
    .A1(\r1.regblock[13][30] ),
    .A2(\r1.regblock[14][30] ),
    .A3(\r1.regblock[15][30] ),
    .S0(net27),
    .S1(net20),
    .X(_01189_));
 sky130_fd_sc_hd__mux4_2 _13666_ (.A0(_01186_),
    .A1(_01187_),
    .A2(_01188_),
    .A3(_01189_),
    .S0(net14),
    .S1(net12),
    .X(_01190_));
 sky130_fd_sc_hd__mux4_1 _13667_ (.A0(\r1.regblock[16][30] ),
    .A1(\r1.regblock[17][30] ),
    .A2(\r1.regblock[18][30] ),
    .A3(\r1.regblock[19][30] ),
    .S0(net28),
    .S1(net20),
    .X(_01191_));
 sky130_fd_sc_hd__mux4_1 _13668_ (.A0(\r1.regblock[20][30] ),
    .A1(\r1.regblock[21][30] ),
    .A2(\r1.regblock[22][30] ),
    .A3(\r1.regblock[23][30] ),
    .S0(net28),
    .S1(net20),
    .X(_01192_));
 sky130_fd_sc_hd__mux4_2 _13669_ (.A0(\r1.regblock[24][30] ),
    .A1(\r1.regblock[25][30] ),
    .A2(\r1.regblock[26][30] ),
    .A3(\r1.regblock[27][30] ),
    .S0(net28),
    .S1(net20),
    .X(_01193_));
 sky130_fd_sc_hd__mux4_2 _13670_ (.A0(\r1.regblock[28][30] ),
    .A1(\r1.regblock[29][30] ),
    .A2(\r1.regblock[30][30] ),
    .A3(\r1.regblock[31][30] ),
    .S0(net28),
    .S1(net20),
    .X(_01194_));
 sky130_fd_sc_hd__mux4_1 _13671_ (.A0(_01191_),
    .A1(_01192_),
    .A2(_01193_),
    .A3(_01194_),
    .S0(net15),
    .S1(\c1.instruction1[18] ),
    .X(_01195_));
 sky130_fd_sc_hd__mux4_1 _13672_ (.A0(\r1.regblock[0][29] ),
    .A1(\r1.regblock[1][29] ),
    .A2(\r1.regblock[2][29] ),
    .A3(\r1.regblock[3][29] ),
    .S0(net27),
    .S1(net19),
    .X(_01174_));
 sky130_fd_sc_hd__mux4_2 _13673_ (.A0(\r1.regblock[4][29] ),
    .A1(\r1.regblock[5][29] ),
    .A2(\r1.regblock[6][29] ),
    .A3(\r1.regblock[7][29] ),
    .S0(net27),
    .S1(net19),
    .X(_01175_));
 sky130_fd_sc_hd__mux4_1 _13674_ (.A0(\r1.regblock[8][29] ),
    .A1(\r1.regblock[9][29] ),
    .A2(\r1.regblock[10][29] ),
    .A3(\r1.regblock[11][29] ),
    .S0(net27),
    .S1(net19),
    .X(_01176_));
 sky130_fd_sc_hd__mux4_1 _13675_ (.A0(\r1.regblock[12][29] ),
    .A1(\r1.regblock[13][29] ),
    .A2(\r1.regblock[14][29] ),
    .A3(\r1.regblock[15][29] ),
    .S0(net27),
    .S1(net19),
    .X(_01177_));
 sky130_fd_sc_hd__mux4_2 _13676_ (.A0(_01174_),
    .A1(_01175_),
    .A2(_01176_),
    .A3(_01177_),
    .S0(net14),
    .S1(net12),
    .X(_01178_));
 sky130_fd_sc_hd__mux4_1 _13677_ (.A0(\r1.regblock[16][29] ),
    .A1(\r1.regblock[17][29] ),
    .A2(\r1.regblock[18][29] ),
    .A3(\r1.regblock[19][29] ),
    .S0(net28),
    .S1(net20),
    .X(_01179_));
 sky130_fd_sc_hd__mux4_2 _13678_ (.A0(\r1.regblock[20][29] ),
    .A1(\r1.regblock[21][29] ),
    .A2(\r1.regblock[22][29] ),
    .A3(\r1.regblock[23][29] ),
    .S0(net28),
    .S1(net20),
    .X(_01180_));
 sky130_fd_sc_hd__mux4_2 _13679_ (.A0(\r1.regblock[24][29] ),
    .A1(\r1.regblock[25][29] ),
    .A2(\r1.regblock[26][29] ),
    .A3(\r1.regblock[27][29] ),
    .S0(net28),
    .S1(net20),
    .X(_01181_));
 sky130_fd_sc_hd__mux4_2 _13680_ (.A0(\r1.regblock[28][29] ),
    .A1(\r1.regblock[29][29] ),
    .A2(\r1.regblock[30][29] ),
    .A3(\r1.regblock[31][29] ),
    .S0(net28),
    .S1(net20),
    .X(_01182_));
 sky130_fd_sc_hd__mux4_1 _13681_ (.A0(_01179_),
    .A1(_01180_),
    .A2(_01181_),
    .A3(_01182_),
    .S0(net15),
    .S1(\c1.instruction1[18] ),
    .X(_01183_));
 sky130_fd_sc_hd__mux4_1 _13682_ (.A0(\r1.regblock[0][28] ),
    .A1(\r1.regblock[1][28] ),
    .A2(\r1.regblock[2][28] ),
    .A3(\r1.regblock[3][28] ),
    .S0(net26),
    .S1(net19),
    .X(_01162_));
 sky130_fd_sc_hd__mux4_2 _13683_ (.A0(\r1.regblock[4][28] ),
    .A1(\r1.regblock[5][28] ),
    .A2(\r1.regblock[6][28] ),
    .A3(\r1.regblock[7][28] ),
    .S0(net26),
    .S1(net19),
    .X(_01163_));
 sky130_fd_sc_hd__mux4_2 _13684_ (.A0(\r1.regblock[8][28] ),
    .A1(\r1.regblock[9][28] ),
    .A2(\r1.regblock[10][28] ),
    .A3(\r1.regblock[11][28] ),
    .S0(net26),
    .S1(net18),
    .X(_01164_));
 sky130_fd_sc_hd__mux4_1 _13685_ (.A0(\r1.regblock[12][28] ),
    .A1(\r1.regblock[13][28] ),
    .A2(\r1.regblock[14][28] ),
    .A3(\r1.regblock[15][28] ),
    .S0(net26),
    .S1(net19),
    .X(_01165_));
 sky130_fd_sc_hd__mux4_2 _13686_ (.A0(_01162_),
    .A1(_01163_),
    .A2(_01164_),
    .A3(_01165_),
    .S0(net14),
    .S1(net12),
    .X(_01166_));
 sky130_fd_sc_hd__mux4_2 _13687_ (.A0(\r1.regblock[16][28] ),
    .A1(\r1.regblock[17][28] ),
    .A2(\r1.regblock[18][28] ),
    .A3(\r1.regblock[19][28] ),
    .S0(net27),
    .S1(net19),
    .X(_01167_));
 sky130_fd_sc_hd__mux4_2 _13688_ (.A0(\r1.regblock[20][28] ),
    .A1(\r1.regblock[21][28] ),
    .A2(\r1.regblock[22][28] ),
    .A3(\r1.regblock[23][28] ),
    .S0(net27),
    .S1(net19),
    .X(_01168_));
 sky130_fd_sc_hd__mux4_2 _13689_ (.A0(\r1.regblock[24][28] ),
    .A1(\r1.regblock[25][28] ),
    .A2(\r1.regblock[26][28] ),
    .A3(\r1.regblock[27][28] ),
    .S0(net27),
    .S1(net19),
    .X(_01169_));
 sky130_fd_sc_hd__mux4_2 _13690_ (.A0(\r1.regblock[28][28] ),
    .A1(\r1.regblock[29][28] ),
    .A2(\r1.regblock[30][28] ),
    .A3(\r1.regblock[31][28] ),
    .S0(net26),
    .S1(net19),
    .X(_01170_));
 sky130_fd_sc_hd__mux4_1 _13691_ (.A0(_01167_),
    .A1(_01168_),
    .A2(_01169_),
    .A3(_01170_),
    .S0(net14),
    .S1(net12),
    .X(_01171_));
 sky130_fd_sc_hd__mux4_1 _13692_ (.A0(\r1.regblock[0][27] ),
    .A1(\r1.regblock[1][27] ),
    .A2(\r1.regblock[2][27] ),
    .A3(\r1.regblock[3][27] ),
    .S0(net26),
    .S1(net19),
    .X(_01150_));
 sky130_fd_sc_hd__mux4_2 _13693_ (.A0(\r1.regblock[4][27] ),
    .A1(\r1.regblock[5][27] ),
    .A2(\r1.regblock[6][27] ),
    .A3(\r1.regblock[7][27] ),
    .S0(net26),
    .S1(net19),
    .X(_01151_));
 sky130_fd_sc_hd__mux4_2 _13694_ (.A0(\r1.regblock[8][27] ),
    .A1(\r1.regblock[9][27] ),
    .A2(\r1.regblock[10][27] ),
    .A3(\r1.regblock[11][27] ),
    .S0(net26),
    .S1(net18),
    .X(_01152_));
 sky130_fd_sc_hd__mux4_2 _13695_ (.A0(\r1.regblock[12][27] ),
    .A1(\r1.regblock[13][27] ),
    .A2(\r1.regblock[14][27] ),
    .A3(\r1.regblock[15][27] ),
    .S0(net26),
    .S1(net19),
    .X(_01153_));
 sky130_fd_sc_hd__mux4_2 _13696_ (.A0(_01150_),
    .A1(_01151_),
    .A2(_01152_),
    .A3(_01153_),
    .S0(net14),
    .S1(net12),
    .X(_01154_));
 sky130_fd_sc_hd__mux4_2 _13697_ (.A0(\r1.regblock[16][27] ),
    .A1(\r1.regblock[17][27] ),
    .A2(\r1.regblock[18][27] ),
    .A3(\r1.regblock[19][27] ),
    .S0(net27),
    .S1(net19),
    .X(_01155_));
 sky130_fd_sc_hd__mux4_1 _13698_ (.A0(\r1.regblock[20][27] ),
    .A1(\r1.regblock[21][27] ),
    .A2(\r1.regblock[22][27] ),
    .A3(\r1.regblock[23][27] ),
    .S0(net27),
    .S1(net19),
    .X(_01156_));
 sky130_fd_sc_hd__mux4_1 _13699_ (.A0(\r1.regblock[24][27] ),
    .A1(\r1.regblock[25][27] ),
    .A2(\r1.regblock[26][27] ),
    .A3(\r1.regblock[27][27] ),
    .S0(net27),
    .S1(net19),
    .X(_01157_));
 sky130_fd_sc_hd__mux4_2 _13700_ (.A0(\r1.regblock[28][27] ),
    .A1(\r1.regblock[29][27] ),
    .A2(\r1.regblock[30][27] ),
    .A3(\r1.regblock[31][27] ),
    .S0(net26),
    .S1(net19),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_1 _13701_ (.A0(_01155_),
    .A1(_01156_),
    .A2(_01157_),
    .A3(_01158_),
    .S0(net14),
    .S1(net12),
    .X(_01159_));
 sky130_fd_sc_hd__mux4_1 _13702_ (.A0(\r1.regblock[0][26] ),
    .A1(\r1.regblock[1][26] ),
    .A2(\r1.regblock[2][26] ),
    .A3(\r1.regblock[3][26] ),
    .S0(net26),
    .S1(net18),
    .X(_01138_));
 sky130_fd_sc_hd__mux4_2 _13703_ (.A0(\r1.regblock[4][26] ),
    .A1(\r1.regblock[5][26] ),
    .A2(\r1.regblock[6][26] ),
    .A3(\r1.regblock[7][26] ),
    .S0(net26),
    .S1(net19),
    .X(_01139_));
 sky130_fd_sc_hd__mux4_2 _13704_ (.A0(\r1.regblock[8][26] ),
    .A1(\r1.regblock[9][26] ),
    .A2(\r1.regblock[10][26] ),
    .A3(\r1.regblock[11][26] ),
    .S0(net26),
    .S1(net18),
    .X(_01140_));
 sky130_fd_sc_hd__mux4_2 _13705_ (.A0(\r1.regblock[12][26] ),
    .A1(\r1.regblock[13][26] ),
    .A2(\r1.regblock[14][26] ),
    .A3(\r1.regblock[15][26] ),
    .S0(net26),
    .S1(net19),
    .X(_01141_));
 sky130_fd_sc_hd__mux4_2 _13706_ (.A0(_01138_),
    .A1(_01139_),
    .A2(_01140_),
    .A3(_01141_),
    .S0(net14),
    .S1(net12),
    .X(_01142_));
 sky130_fd_sc_hd__mux4_1 _13707_ (.A0(\r1.regblock[16][26] ),
    .A1(\r1.regblock[17][26] ),
    .A2(\r1.regblock[18][26] ),
    .A3(\r1.regblock[19][26] ),
    .S0(net27),
    .S1(net19),
    .X(_01143_));
 sky130_fd_sc_hd__mux4_2 _13708_ (.A0(\r1.regblock[20][26] ),
    .A1(\r1.regblock[21][26] ),
    .A2(\r1.regblock[22][26] ),
    .A3(\r1.regblock[23][26] ),
    .S0(net27),
    .S1(net19),
    .X(_01144_));
 sky130_fd_sc_hd__mux4_2 _13709_ (.A0(\r1.regblock[24][26] ),
    .A1(\r1.regblock[25][26] ),
    .A2(\r1.regblock[26][26] ),
    .A3(\r1.regblock[27][26] ),
    .S0(net27),
    .S1(net19),
    .X(_01145_));
 sky130_fd_sc_hd__mux4_2 _13710_ (.A0(\r1.regblock[28][26] ),
    .A1(\r1.regblock[29][26] ),
    .A2(\r1.regblock[30][26] ),
    .A3(\r1.regblock[31][26] ),
    .S0(net26),
    .S1(net19),
    .X(_01146_));
 sky130_fd_sc_hd__mux4_1 _13711_ (.A0(_01143_),
    .A1(_01144_),
    .A2(_01145_),
    .A3(_01146_),
    .S0(net14),
    .S1(net12),
    .X(_01147_));
 sky130_fd_sc_hd__mux4_1 _13712_ (.A0(\r1.regblock[0][25] ),
    .A1(\r1.regblock[1][25] ),
    .A2(\r1.regblock[2][25] ),
    .A3(\r1.regblock[3][25] ),
    .S0(net26),
    .S1(net18),
    .X(_01126_));
 sky130_fd_sc_hd__mux4_1 _13713_ (.A0(\r1.regblock[4][25] ),
    .A1(\r1.regblock[5][25] ),
    .A2(\r1.regblock[6][25] ),
    .A3(\r1.regblock[7][25] ),
    .S0(net26),
    .S1(net18),
    .X(_01127_));
 sky130_fd_sc_hd__mux4_2 _13714_ (.A0(\r1.regblock[8][25] ),
    .A1(\r1.regblock[9][25] ),
    .A2(\r1.regblock[10][25] ),
    .A3(\r1.regblock[11][25] ),
    .S0(net26),
    .S1(net18),
    .X(_01128_));
 sky130_fd_sc_hd__mux4_2 _13715_ (.A0(\r1.regblock[12][25] ),
    .A1(\r1.regblock[13][25] ),
    .A2(\r1.regblock[14][25] ),
    .A3(\r1.regblock[15][25] ),
    .S0(net26),
    .S1(net18),
    .X(_01129_));
 sky130_fd_sc_hd__mux4_2 _13716_ (.A0(_01126_),
    .A1(_01127_),
    .A2(_01128_),
    .A3(_01129_),
    .S0(net14),
    .S1(net12),
    .X(_01130_));
 sky130_fd_sc_hd__mux4_2 _13717_ (.A0(\r1.regblock[16][25] ),
    .A1(\r1.regblock[17][25] ),
    .A2(\r1.regblock[18][25] ),
    .A3(\r1.regblock[19][25] ),
    .S0(net26),
    .S1(net19),
    .X(_01131_));
 sky130_fd_sc_hd__mux4_1 _13718_ (.A0(\r1.regblock[20][25] ),
    .A1(\r1.regblock[21][25] ),
    .A2(\r1.regblock[22][25] ),
    .A3(\r1.regblock[23][25] ),
    .S0(net26),
    .S1(net19),
    .X(_01132_));
 sky130_fd_sc_hd__mux4_2 _13719_ (.A0(\r1.regblock[24][25] ),
    .A1(\r1.regblock[25][25] ),
    .A2(\r1.regblock[26][25] ),
    .A3(\r1.regblock[27][25] ),
    .S0(net27),
    .S1(net19),
    .X(_01133_));
 sky130_fd_sc_hd__mux4_2 _13720_ (.A0(\r1.regblock[28][25] ),
    .A1(\r1.regblock[29][25] ),
    .A2(\r1.regblock[30][25] ),
    .A3(\r1.regblock[31][25] ),
    .S0(net27),
    .S1(net19),
    .X(_01134_));
 sky130_fd_sc_hd__mux4_1 _13721_ (.A0(_01131_),
    .A1(_01132_),
    .A2(_01133_),
    .A3(_01134_),
    .S0(net14),
    .S1(net12),
    .X(_01135_));
 sky130_fd_sc_hd__mux4_1 _13722_ (.A0(\r1.regblock[0][24] ),
    .A1(\r1.regblock[1][24] ),
    .A2(\r1.regblock[2][24] ),
    .A3(\r1.regblock[3][24] ),
    .S0(net26),
    .S1(net18),
    .X(_01114_));
 sky130_fd_sc_hd__mux4_2 _13723_ (.A0(\r1.regblock[4][24] ),
    .A1(\r1.regblock[5][24] ),
    .A2(\r1.regblock[6][24] ),
    .A3(\r1.regblock[7][24] ),
    .S0(net26),
    .S1(net18),
    .X(_01115_));
 sky130_fd_sc_hd__mux4_2 _13724_ (.A0(\r1.regblock[8][24] ),
    .A1(\r1.regblock[9][24] ),
    .A2(\r1.regblock[10][24] ),
    .A3(\r1.regblock[11][24] ),
    .S0(net25),
    .S1(net18),
    .X(_01116_));
 sky130_fd_sc_hd__mux4_1 _13725_ (.A0(\r1.regblock[12][24] ),
    .A1(\r1.regblock[13][24] ),
    .A2(\r1.regblock[14][24] ),
    .A3(\r1.regblock[15][24] ),
    .S0(net26),
    .S1(net18),
    .X(_01117_));
 sky130_fd_sc_hd__mux4_2 _13726_ (.A0(_01114_),
    .A1(_01115_),
    .A2(_01116_),
    .A3(_01117_),
    .S0(net14),
    .S1(net12),
    .X(_01118_));
 sky130_fd_sc_hd__mux4_2 _13727_ (.A0(\r1.regblock[16][24] ),
    .A1(\r1.regblock[17][24] ),
    .A2(\r1.regblock[18][24] ),
    .A3(\r1.regblock[19][24] ),
    .S0(net26),
    .S1(net19),
    .X(_01119_));
 sky130_fd_sc_hd__mux4_2 _13728_ (.A0(\r1.regblock[20][24] ),
    .A1(\r1.regblock[21][24] ),
    .A2(\r1.regblock[22][24] ),
    .A3(\r1.regblock[23][24] ),
    .S0(net27),
    .S1(net19),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_1 _13729_ (.A0(\r1.regblock[24][24] ),
    .A1(\r1.regblock[25][24] ),
    .A2(\r1.regblock[26][24] ),
    .A3(\r1.regblock[27][24] ),
    .S0(net27),
    .S1(net19),
    .X(_01121_));
 sky130_fd_sc_hd__mux4_1 _13730_ (.A0(\r1.regblock[28][24] ),
    .A1(\r1.regblock[29][24] ),
    .A2(\r1.regblock[30][24] ),
    .A3(\r1.regblock[31][24] ),
    .S0(net27),
    .S1(net19),
    .X(_01122_));
 sky130_fd_sc_hd__mux4_1 _13731_ (.A0(_01119_),
    .A1(_01120_),
    .A2(_01121_),
    .A3(_01122_),
    .S0(net14),
    .S1(net12),
    .X(_01123_));
 sky130_fd_sc_hd__mux4_1 _13732_ (.A0(\r1.regblock[0][23] ),
    .A1(\r1.regblock[1][23] ),
    .A2(\r1.regblock[2][23] ),
    .A3(\r1.regblock[3][23] ),
    .S0(net26),
    .S1(net18),
    .X(_01102_));
 sky130_fd_sc_hd__mux4_2 _13733_ (.A0(\r1.regblock[4][23] ),
    .A1(\r1.regblock[5][23] ),
    .A2(\r1.regblock[6][23] ),
    .A3(\r1.regblock[7][23] ),
    .S0(net26),
    .S1(net18),
    .X(_01103_));
 sky130_fd_sc_hd__mux4_2 _13734_ (.A0(\r1.regblock[8][23] ),
    .A1(\r1.regblock[9][23] ),
    .A2(\r1.regblock[10][23] ),
    .A3(\r1.regblock[11][23] ),
    .S0(net25),
    .S1(net18),
    .X(_01104_));
 sky130_fd_sc_hd__mux4_1 _13735_ (.A0(\r1.regblock[12][23] ),
    .A1(\r1.regblock[13][23] ),
    .A2(\r1.regblock[14][23] ),
    .A3(\r1.regblock[15][23] ),
    .S0(net26),
    .S1(net18),
    .X(_01105_));
 sky130_fd_sc_hd__mux4_2 _13736_ (.A0(_01102_),
    .A1(_01103_),
    .A2(_01104_),
    .A3(_01105_),
    .S0(net14),
    .S1(net12),
    .X(_01106_));
 sky130_fd_sc_hd__mux4_2 _13737_ (.A0(\r1.regblock[16][23] ),
    .A1(\r1.regblock[17][23] ),
    .A2(\r1.regblock[18][23] ),
    .A3(\r1.regblock[19][23] ),
    .S0(net26),
    .S1(net19),
    .X(_01107_));
 sky130_fd_sc_hd__mux4_1 _13738_ (.A0(\r1.regblock[20][23] ),
    .A1(\r1.regblock[21][23] ),
    .A2(\r1.regblock[22][23] ),
    .A3(\r1.regblock[23][23] ),
    .S0(net27),
    .S1(net19),
    .X(_01108_));
 sky130_fd_sc_hd__mux4_2 _13739_ (.A0(\r1.regblock[24][23] ),
    .A1(\r1.regblock[25][23] ),
    .A2(\r1.regblock[26][23] ),
    .A3(\r1.regblock[27][23] ),
    .S0(net27),
    .S1(net19),
    .X(_01109_));
 sky130_fd_sc_hd__mux4_2 _13740_ (.A0(\r1.regblock[28][23] ),
    .A1(\r1.regblock[29][23] ),
    .A2(\r1.regblock[30][23] ),
    .A3(\r1.regblock[31][23] ),
    .S0(net27),
    .S1(net19),
    .X(_01110_));
 sky130_fd_sc_hd__mux4_1 _13741_ (.A0(_01107_),
    .A1(_01108_),
    .A2(_01109_),
    .A3(_01110_),
    .S0(net14),
    .S1(net12),
    .X(_01111_));
 sky130_fd_sc_hd__mux4_1 _13742_ (.A0(\r1.regblock[0][22] ),
    .A1(\r1.regblock[1][22] ),
    .A2(\r1.regblock[2][22] ),
    .A3(\r1.regblock[3][22] ),
    .S0(net25),
    .S1(net18),
    .X(_01090_));
 sky130_fd_sc_hd__mux4_2 _13743_ (.A0(\r1.regblock[4][22] ),
    .A1(\r1.regblock[5][22] ),
    .A2(\r1.regblock[6][22] ),
    .A3(\r1.regblock[7][22] ),
    .S0(net25),
    .S1(net18),
    .X(_01091_));
 sky130_fd_sc_hd__mux4_2 _13744_ (.A0(\r1.regblock[8][22] ),
    .A1(\r1.regblock[9][22] ),
    .A2(\r1.regblock[10][22] ),
    .A3(\r1.regblock[11][22] ),
    .S0(net25),
    .S1(net18),
    .X(_01092_));
 sky130_fd_sc_hd__mux4_1 _13745_ (.A0(\r1.regblock[12][22] ),
    .A1(\r1.regblock[13][22] ),
    .A2(\r1.regblock[14][22] ),
    .A3(\r1.regblock[15][22] ),
    .S0(net25),
    .S1(net18),
    .X(_01093_));
 sky130_fd_sc_hd__mux4_2 _13746_ (.A0(_01090_),
    .A1(_01091_),
    .A2(_01092_),
    .A3(_01093_),
    .S0(net14),
    .S1(net12),
    .X(_01094_));
 sky130_fd_sc_hd__mux4_2 _13747_ (.A0(\r1.regblock[16][22] ),
    .A1(\r1.regblock[17][22] ),
    .A2(\r1.regblock[18][22] ),
    .A3(\r1.regblock[19][22] ),
    .S0(net25),
    .S1(net18),
    .X(_01095_));
 sky130_fd_sc_hd__mux4_2 _13748_ (.A0(\r1.regblock[20][22] ),
    .A1(\r1.regblock[21][22] ),
    .A2(\r1.regblock[22][22] ),
    .A3(\r1.regblock[23][22] ),
    .S0(net25),
    .S1(net18),
    .X(_01096_));
 sky130_fd_sc_hd__mux4_2 _13749_ (.A0(\r1.regblock[24][22] ),
    .A1(\r1.regblock[25][22] ),
    .A2(\r1.regblock[26][22] ),
    .A3(\r1.regblock[27][22] ),
    .S0(net25),
    .S1(net18),
    .X(_01097_));
 sky130_fd_sc_hd__mux4_1 _13750_ (.A0(\r1.regblock[28][22] ),
    .A1(\r1.regblock[29][22] ),
    .A2(\r1.regblock[30][22] ),
    .A3(\r1.regblock[31][22] ),
    .S0(net25),
    .S1(net18),
    .X(_01098_));
 sky130_fd_sc_hd__mux4_1 _13751_ (.A0(_01095_),
    .A1(_01096_),
    .A2(_01097_),
    .A3(_01098_),
    .S0(net14),
    .S1(net12),
    .X(_01099_));
 sky130_fd_sc_hd__mux4_1 _13752_ (.A0(\r1.regblock[0][21] ),
    .A1(\r1.regblock[1][21] ),
    .A2(\r1.regblock[2][21] ),
    .A3(\r1.regblock[3][21] ),
    .S0(net25),
    .S1(net18),
    .X(_01078_));
 sky130_fd_sc_hd__mux4_2 _13753_ (.A0(\r1.regblock[4][21] ),
    .A1(\r1.regblock[5][21] ),
    .A2(\r1.regblock[6][21] ),
    .A3(\r1.regblock[7][21] ),
    .S0(net25),
    .S1(net18),
    .X(_01079_));
 sky130_fd_sc_hd__mux4_2 _13754_ (.A0(\r1.regblock[8][21] ),
    .A1(\r1.regblock[9][21] ),
    .A2(\r1.regblock[10][21] ),
    .A3(\r1.regblock[11][21] ),
    .S0(net25),
    .S1(net18),
    .X(_01080_));
 sky130_fd_sc_hd__mux4_1 _13755_ (.A0(\r1.regblock[12][21] ),
    .A1(\r1.regblock[13][21] ),
    .A2(\r1.regblock[14][21] ),
    .A3(\r1.regblock[15][21] ),
    .S0(net25),
    .S1(net18),
    .X(_01081_));
 sky130_fd_sc_hd__mux4_2 _13756_ (.A0(_01078_),
    .A1(_01079_),
    .A2(_01080_),
    .A3(_01081_),
    .S0(net14),
    .S1(net12),
    .X(_01082_));
 sky130_fd_sc_hd__mux4_2 _13757_ (.A0(\r1.regblock[16][21] ),
    .A1(\r1.regblock[17][21] ),
    .A2(\r1.regblock[18][21] ),
    .A3(\r1.regblock[19][21] ),
    .S0(net25),
    .S1(net18),
    .X(_01083_));
 sky130_fd_sc_hd__mux4_1 _13758_ (.A0(\r1.regblock[20][21] ),
    .A1(\r1.regblock[21][21] ),
    .A2(\r1.regblock[22][21] ),
    .A3(\r1.regblock[23][21] ),
    .S0(net25),
    .S1(net18),
    .X(_01084_));
 sky130_fd_sc_hd__mux4_2 _13759_ (.A0(\r1.regblock[24][21] ),
    .A1(\r1.regblock[25][21] ),
    .A2(\r1.regblock[26][21] ),
    .A3(\r1.regblock[27][21] ),
    .S0(net25),
    .S1(net18),
    .X(_01085_));
 sky130_fd_sc_hd__mux4_1 _13760_ (.A0(\r1.regblock[28][21] ),
    .A1(\r1.regblock[29][21] ),
    .A2(\r1.regblock[30][21] ),
    .A3(\r1.regblock[31][21] ),
    .S0(net25),
    .S1(net18),
    .X(_01086_));
 sky130_fd_sc_hd__mux4_1 _13761_ (.A0(_01083_),
    .A1(_01084_),
    .A2(_01085_),
    .A3(_01086_),
    .S0(net14),
    .S1(net12),
    .X(_01087_));
 sky130_fd_sc_hd__mux4_1 _13762_ (.A0(\r1.regblock[0][20] ),
    .A1(\r1.regblock[1][20] ),
    .A2(\r1.regblock[2][20] ),
    .A3(\r1.regblock[3][20] ),
    .S0(net25),
    .S1(net18),
    .X(_01066_));
 sky130_fd_sc_hd__mux4_2 _13763_ (.A0(\r1.regblock[4][20] ),
    .A1(\r1.regblock[5][20] ),
    .A2(\r1.regblock[6][20] ),
    .A3(\r1.regblock[7][20] ),
    .S0(net25),
    .S1(net18),
    .X(_01067_));
 sky130_fd_sc_hd__mux4_1 _13764_ (.A0(\r1.regblock[8][20] ),
    .A1(\r1.regblock[9][20] ),
    .A2(\r1.regblock[10][20] ),
    .A3(\r1.regblock[11][20] ),
    .S0(net25),
    .S1(net18),
    .X(_01068_));
 sky130_fd_sc_hd__mux4_2 _13765_ (.A0(\r1.regblock[12][20] ),
    .A1(\r1.regblock[13][20] ),
    .A2(\r1.regblock[14][20] ),
    .A3(\r1.regblock[15][20] ),
    .S0(net25),
    .S1(net18),
    .X(_01069_));
 sky130_fd_sc_hd__mux4_2 _13766_ (.A0(_01066_),
    .A1(_01067_),
    .A2(_01068_),
    .A3(_01069_),
    .S0(net14),
    .S1(net12),
    .X(_01070_));
 sky130_fd_sc_hd__mux4_2 _13767_ (.A0(\r1.regblock[16][20] ),
    .A1(\r1.regblock[17][20] ),
    .A2(\r1.regblock[18][20] ),
    .A3(\r1.regblock[19][20] ),
    .S0(net25),
    .S1(net18),
    .X(_01071_));
 sky130_fd_sc_hd__mux4_2 _13768_ (.A0(\r1.regblock[20][20] ),
    .A1(\r1.regblock[21][20] ),
    .A2(\r1.regblock[22][20] ),
    .A3(\r1.regblock[23][20] ),
    .S0(net25),
    .S1(net18),
    .X(_01072_));
 sky130_fd_sc_hd__mux4_1 _13769_ (.A0(\r1.regblock[24][20] ),
    .A1(\r1.regblock[25][20] ),
    .A2(\r1.regblock[26][20] ),
    .A3(\r1.regblock[27][20] ),
    .S0(net25),
    .S1(net18),
    .X(_01073_));
 sky130_fd_sc_hd__mux4_1 _13770_ (.A0(\r1.regblock[28][20] ),
    .A1(\r1.regblock[29][20] ),
    .A2(\r1.regblock[30][20] ),
    .A3(\r1.regblock[31][20] ),
    .S0(net25),
    .S1(net18),
    .X(_01074_));
 sky130_fd_sc_hd__mux4_1 _13771_ (.A0(_01071_),
    .A1(_01072_),
    .A2(_01073_),
    .A3(_01074_),
    .S0(net14),
    .S1(net12),
    .X(_01075_));
 sky130_fd_sc_hd__mux4_1 _13772_ (.A0(\r1.regblock[0][19] ),
    .A1(\r1.regblock[1][19] ),
    .A2(\r1.regblock[2][19] ),
    .A3(\r1.regblock[3][19] ),
    .S0(net23),
    .S1(net17),
    .X(_01054_));
 sky130_fd_sc_hd__mux4_2 _13773_ (.A0(\r1.regblock[4][19] ),
    .A1(\r1.regblock[5][19] ),
    .A2(\r1.regblock[6][19] ),
    .A3(\r1.regblock[7][19] ),
    .S0(net24),
    .S1(net16),
    .X(_01055_));
 sky130_fd_sc_hd__mux4_1 _13774_ (.A0(\r1.regblock[8][19] ),
    .A1(\r1.regblock[9][19] ),
    .A2(\r1.regblock[10][19] ),
    .A3(\r1.regblock[11][19] ),
    .S0(net24),
    .S1(net17),
    .X(_01056_));
 sky130_fd_sc_hd__mux4_1 _13775_ (.A0(\r1.regblock[12][19] ),
    .A1(\r1.regblock[13][19] ),
    .A2(\r1.regblock[14][19] ),
    .A3(\r1.regblock[15][19] ),
    .S0(net23),
    .S1(net17),
    .X(_01057_));
 sky130_fd_sc_hd__mux4_2 _13776_ (.A0(_01054_),
    .A1(_01055_),
    .A2(_01056_),
    .A3(_01057_),
    .S0(net15),
    .S1(net13),
    .X(_01058_));
 sky130_fd_sc_hd__mux4_2 _13777_ (.A0(\r1.regblock[16][19] ),
    .A1(\r1.regblock[17][19] ),
    .A2(\r1.regblock[18][19] ),
    .A3(\r1.regblock[19][19] ),
    .S0(net23),
    .S1(net17),
    .X(_01059_));
 sky130_fd_sc_hd__mux4_1 _13778_ (.A0(\r1.regblock[20][19] ),
    .A1(\r1.regblock[21][19] ),
    .A2(\r1.regblock[22][19] ),
    .A3(\r1.regblock[23][19] ),
    .S0(net23),
    .S1(net17),
    .X(_01060_));
 sky130_fd_sc_hd__mux4_2 _13779_ (.A0(\r1.regblock[24][19] ),
    .A1(\r1.regblock[25][19] ),
    .A2(\r1.regblock[26][19] ),
    .A3(\r1.regblock[27][19] ),
    .S0(net23),
    .S1(net17),
    .X(_01061_));
 sky130_fd_sc_hd__mux4_2 _13780_ (.A0(\r1.regblock[28][19] ),
    .A1(\r1.regblock[29][19] ),
    .A2(\r1.regblock[30][19] ),
    .A3(\r1.regblock[31][19] ),
    .S0(net23),
    .S1(net17),
    .X(_01062_));
 sky130_fd_sc_hd__mux4_1 _13781_ (.A0(_01059_),
    .A1(_01060_),
    .A2(_01061_),
    .A3(_01062_),
    .S0(net15),
    .S1(\c1.instruction1[18] ),
    .X(_01063_));
 sky130_fd_sc_hd__mux4_1 _13782_ (.A0(\r1.regblock[0][18] ),
    .A1(\r1.regblock[1][18] ),
    .A2(\r1.regblock[2][18] ),
    .A3(\r1.regblock[3][18] ),
    .S0(net23),
    .S1(net17),
    .X(_01042_));
 sky130_fd_sc_hd__mux4_2 _13783_ (.A0(\r1.regblock[4][18] ),
    .A1(\r1.regblock[5][18] ),
    .A2(\r1.regblock[6][18] ),
    .A3(\r1.regblock[7][18] ),
    .S0(net24),
    .S1(net16),
    .X(_01043_));
 sky130_fd_sc_hd__mux4_1 _13784_ (.A0(\r1.regblock[8][18] ),
    .A1(\r1.regblock[9][18] ),
    .A2(\r1.regblock[10][18] ),
    .A3(\r1.regblock[11][18] ),
    .S0(net23),
    .S1(net17),
    .X(_01044_));
 sky130_fd_sc_hd__mux4_1 _13785_ (.A0(\r1.regblock[12][18] ),
    .A1(\r1.regblock[13][18] ),
    .A2(\r1.regblock[14][18] ),
    .A3(\r1.regblock[15][18] ),
    .S0(net23),
    .S1(net17),
    .X(_01045_));
 sky130_fd_sc_hd__mux4_2 _13786_ (.A0(_01042_),
    .A1(_01043_),
    .A2(_01044_),
    .A3(_01045_),
    .S0(net15),
    .S1(net13),
    .X(_01046_));
 sky130_fd_sc_hd__mux4_2 _13787_ (.A0(\r1.regblock[16][18] ),
    .A1(\r1.regblock[17][18] ),
    .A2(\r1.regblock[18][18] ),
    .A3(\r1.regblock[19][18] ),
    .S0(net23),
    .S1(net17),
    .X(_01047_));
 sky130_fd_sc_hd__mux4_1 _13788_ (.A0(\r1.regblock[20][18] ),
    .A1(\r1.regblock[21][18] ),
    .A2(\r1.regblock[22][18] ),
    .A3(\r1.regblock[23][18] ),
    .S0(net23),
    .S1(net17),
    .X(_01048_));
 sky130_fd_sc_hd__mux4_2 _13789_ (.A0(\r1.regblock[24][18] ),
    .A1(\r1.regblock[25][18] ),
    .A2(\r1.regblock[26][18] ),
    .A3(\r1.regblock[27][18] ),
    .S0(net23),
    .S1(net17),
    .X(_01049_));
 sky130_fd_sc_hd__mux4_2 _13790_ (.A0(\r1.regblock[28][18] ),
    .A1(\r1.regblock[29][18] ),
    .A2(\r1.regblock[30][18] ),
    .A3(\r1.regblock[31][18] ),
    .S0(net23),
    .S1(net17),
    .X(_01050_));
 sky130_fd_sc_hd__mux4_1 _13791_ (.A0(_01047_),
    .A1(_01048_),
    .A2(_01049_),
    .A3(_01050_),
    .S0(net15),
    .S1(net13),
    .X(_01051_));
 sky130_fd_sc_hd__mux4_1 _13792_ (.A0(\r1.regblock[0][17] ),
    .A1(\r1.regblock[1][17] ),
    .A2(\r1.regblock[2][17] ),
    .A3(\r1.regblock[3][17] ),
    .S0(net23),
    .S1(net17),
    .X(_01030_));
 sky130_fd_sc_hd__mux4_2 _13793_ (.A0(\r1.regblock[4][17] ),
    .A1(\r1.regblock[5][17] ),
    .A2(\r1.regblock[6][17] ),
    .A3(\r1.regblock[7][17] ),
    .S0(net24),
    .S1(net16),
    .X(_01031_));
 sky130_fd_sc_hd__mux4_1 _13794_ (.A0(\r1.regblock[8][17] ),
    .A1(\r1.regblock[9][17] ),
    .A2(\r1.regblock[10][17] ),
    .A3(\r1.regblock[11][17] ),
    .S0(net23),
    .S1(net17),
    .X(_01032_));
 sky130_fd_sc_hd__mux4_1 _13795_ (.A0(\r1.regblock[12][17] ),
    .A1(\r1.regblock[13][17] ),
    .A2(\r1.regblock[14][17] ),
    .A3(\r1.regblock[15][17] ),
    .S0(net23),
    .S1(net17),
    .X(_01033_));
 sky130_fd_sc_hd__mux4_2 _13796_ (.A0(_01030_),
    .A1(_01031_),
    .A2(_01032_),
    .A3(_01033_),
    .S0(net15),
    .S1(net13),
    .X(_01034_));
 sky130_fd_sc_hd__mux4_2 _13797_ (.A0(\r1.regblock[16][17] ),
    .A1(\r1.regblock[17][17] ),
    .A2(\r1.regblock[18][17] ),
    .A3(\r1.regblock[19][17] ),
    .S0(net23),
    .S1(net17),
    .X(_01035_));
 sky130_fd_sc_hd__mux4_1 _13798_ (.A0(\r1.regblock[20][17] ),
    .A1(\r1.regblock[21][17] ),
    .A2(\r1.regblock[22][17] ),
    .A3(\r1.regblock[23][17] ),
    .S0(net23),
    .S1(net17),
    .X(_01036_));
 sky130_fd_sc_hd__mux4_2 _13799_ (.A0(\r1.regblock[24][17] ),
    .A1(\r1.regblock[25][17] ),
    .A2(\r1.regblock[26][17] ),
    .A3(\r1.regblock[27][17] ),
    .S0(net23),
    .S1(net17),
    .X(_01037_));
 sky130_fd_sc_hd__mux4_2 _13800_ (.A0(\r1.regblock[28][17] ),
    .A1(\r1.regblock[29][17] ),
    .A2(\r1.regblock[30][17] ),
    .A3(\r1.regblock[31][17] ),
    .S0(net23),
    .S1(net17),
    .X(_01038_));
 sky130_fd_sc_hd__mux4_1 _13801_ (.A0(_01035_),
    .A1(_01036_),
    .A2(_01037_),
    .A3(_01038_),
    .S0(net15),
    .S1(net13),
    .X(_01039_));
 sky130_fd_sc_hd__mux4_2 _13802_ (.A0(\r1.regblock[0][16] ),
    .A1(\r1.regblock[1][16] ),
    .A2(\r1.regblock[2][16] ),
    .A3(\r1.regblock[3][16] ),
    .S0(net23),
    .S1(net17),
    .X(_01018_));
 sky130_fd_sc_hd__mux4_2 _13803_ (.A0(\r1.regblock[4][16] ),
    .A1(\r1.regblock[5][16] ),
    .A2(\r1.regblock[6][16] ),
    .A3(\r1.regblock[7][16] ),
    .S0(net24),
    .S1(net16),
    .X(_01019_));
 sky130_fd_sc_hd__mux4_1 _13804_ (.A0(\r1.regblock[8][16] ),
    .A1(\r1.regblock[9][16] ),
    .A2(\r1.regblock[10][16] ),
    .A3(\r1.regblock[11][16] ),
    .S0(net23),
    .S1(net17),
    .X(_01020_));
 sky130_fd_sc_hd__mux4_1 _13805_ (.A0(\r1.regblock[12][16] ),
    .A1(\r1.regblock[13][16] ),
    .A2(\r1.regblock[14][16] ),
    .A3(\r1.regblock[15][16] ),
    .S0(net23),
    .S1(net17),
    .X(_01021_));
 sky130_fd_sc_hd__mux4_2 _13806_ (.A0(_01018_),
    .A1(_01019_),
    .A2(_01020_),
    .A3(_01021_),
    .S0(net15),
    .S1(net13),
    .X(_01022_));
 sky130_fd_sc_hd__mux4_2 _13807_ (.A0(\r1.regblock[16][16] ),
    .A1(\r1.regblock[17][16] ),
    .A2(\r1.regblock[18][16] ),
    .A3(\r1.regblock[19][16] ),
    .S0(net22),
    .S1(net16),
    .X(_01023_));
 sky130_fd_sc_hd__mux4_2 _13808_ (.A0(\r1.regblock[20][16] ),
    .A1(\r1.regblock[21][16] ),
    .A2(\r1.regblock[22][16] ),
    .A3(\r1.regblock[23][16] ),
    .S0(net22),
    .S1(net16),
    .X(_01024_));
 sky130_fd_sc_hd__mux4_2 _13809_ (.A0(\r1.regblock[24][16] ),
    .A1(\r1.regblock[25][16] ),
    .A2(\r1.regblock[26][16] ),
    .A3(\r1.regblock[27][16] ),
    .S0(net22),
    .S1(net16),
    .X(_01025_));
 sky130_fd_sc_hd__mux4_1 _13810_ (.A0(\r1.regblock[28][16] ),
    .A1(\r1.regblock[29][16] ),
    .A2(\r1.regblock[30][16] ),
    .A3(\r1.regblock[31][16] ),
    .S0(net22),
    .S1(net16),
    .X(_01026_));
 sky130_fd_sc_hd__mux4_2 _13811_ (.A0(_01023_),
    .A1(_01024_),
    .A2(_01025_),
    .A3(_01026_),
    .S0(net15),
    .S1(net13),
    .X(_01027_));
 sky130_fd_sc_hd__mux4_1 _13812_ (.A0(\r1.regblock[0][15] ),
    .A1(\r1.regblock[1][15] ),
    .A2(\r1.regblock[2][15] ),
    .A3(\r1.regblock[3][15] ),
    .S0(net23),
    .S1(net17),
    .X(_01006_));
 sky130_fd_sc_hd__mux4_2 _13813_ (.A0(\r1.regblock[4][15] ),
    .A1(\r1.regblock[5][15] ),
    .A2(\r1.regblock[6][15] ),
    .A3(\r1.regblock[7][15] ),
    .S0(net24),
    .S1(net16),
    .X(_01007_));
 sky130_fd_sc_hd__mux4_1 _13814_ (.A0(\r1.regblock[8][15] ),
    .A1(\r1.regblock[9][15] ),
    .A2(\r1.regblock[10][15] ),
    .A3(\r1.regblock[11][15] ),
    .S0(net23),
    .S1(net17),
    .X(_01008_));
 sky130_fd_sc_hd__mux4_2 _13815_ (.A0(\r1.regblock[12][15] ),
    .A1(\r1.regblock[13][15] ),
    .A2(\r1.regblock[14][15] ),
    .A3(\r1.regblock[15][15] ),
    .S0(net23),
    .S1(net17),
    .X(_01009_));
 sky130_fd_sc_hd__mux4_2 _13816_ (.A0(_01006_),
    .A1(_01007_),
    .A2(_01008_),
    .A3(_01009_),
    .S0(net15),
    .S1(net13),
    .X(_01010_));
 sky130_fd_sc_hd__mux4_1 _13817_ (.A0(\r1.regblock[16][15] ),
    .A1(\r1.regblock[17][15] ),
    .A2(\r1.regblock[18][15] ),
    .A3(\r1.regblock[19][15] ),
    .S0(net22),
    .S1(net16),
    .X(_01011_));
 sky130_fd_sc_hd__mux4_2 _13818_ (.A0(\r1.regblock[20][15] ),
    .A1(\r1.regblock[21][15] ),
    .A2(\r1.regblock[22][15] ),
    .A3(\r1.regblock[23][15] ),
    .S0(net22),
    .S1(net16),
    .X(_01012_));
 sky130_fd_sc_hd__mux4_2 _13819_ (.A0(\r1.regblock[24][15] ),
    .A1(\r1.regblock[25][15] ),
    .A2(\r1.regblock[26][15] ),
    .A3(\r1.regblock[27][15] ),
    .S0(net22),
    .S1(net16),
    .X(_01013_));
 sky130_fd_sc_hd__mux4_1 _13820_ (.A0(\r1.regblock[28][15] ),
    .A1(\r1.regblock[29][15] ),
    .A2(\r1.regblock[30][15] ),
    .A3(\r1.regblock[31][15] ),
    .S0(net22),
    .S1(net16),
    .X(_01014_));
 sky130_fd_sc_hd__mux4_1 _13821_ (.A0(_01011_),
    .A1(_01012_),
    .A2(_01013_),
    .A3(_01014_),
    .S0(net15),
    .S1(net13),
    .X(_01015_));
 sky130_fd_sc_hd__mux4_1 _13822_ (.A0(\r1.regblock[0][14] ),
    .A1(\r1.regblock[1][14] ),
    .A2(\r1.regblock[2][14] ),
    .A3(\r1.regblock[3][14] ),
    .S0(net23),
    .S1(net17),
    .X(_00994_));
 sky130_fd_sc_hd__mux4_2 _13823_ (.A0(\r1.regblock[4][14] ),
    .A1(\r1.regblock[5][14] ),
    .A2(\r1.regblock[6][14] ),
    .A3(\r1.regblock[7][14] ),
    .S0(net24),
    .S1(net16),
    .X(_00995_));
 sky130_fd_sc_hd__mux4_1 _13824_ (.A0(\r1.regblock[8][14] ),
    .A1(\r1.regblock[9][14] ),
    .A2(\r1.regblock[10][14] ),
    .A3(\r1.regblock[11][14] ),
    .S0(net23),
    .S1(net17),
    .X(_00996_));
 sky130_fd_sc_hd__mux4_2 _13825_ (.A0(\r1.regblock[12][14] ),
    .A1(\r1.regblock[13][14] ),
    .A2(\r1.regblock[14][14] ),
    .A3(\r1.regblock[15][14] ),
    .S0(net23),
    .S1(net17),
    .X(_00997_));
 sky130_fd_sc_hd__mux4_2 _13826_ (.A0(_00994_),
    .A1(_00995_),
    .A2(_00996_),
    .A3(_00997_),
    .S0(net15),
    .S1(net13),
    .X(_00998_));
 sky130_fd_sc_hd__mux4_1 _13827_ (.A0(\r1.regblock[16][14] ),
    .A1(\r1.regblock[17][14] ),
    .A2(\r1.regblock[18][14] ),
    .A3(\r1.regblock[19][14] ),
    .S0(net22),
    .S1(net16),
    .X(_00999_));
 sky130_fd_sc_hd__mux4_2 _13828_ (.A0(\r1.regblock[20][14] ),
    .A1(\r1.regblock[21][14] ),
    .A2(\r1.regblock[22][14] ),
    .A3(\r1.regblock[23][14] ),
    .S0(net22),
    .S1(net16),
    .X(_01000_));
 sky130_fd_sc_hd__mux4_1 _13829_ (.A0(\r1.regblock[24][14] ),
    .A1(\r1.regblock[25][14] ),
    .A2(\r1.regblock[26][14] ),
    .A3(\r1.regblock[27][14] ),
    .S0(net22),
    .S1(net16),
    .X(_01001_));
 sky130_fd_sc_hd__mux4_1 _13830_ (.A0(\r1.regblock[28][14] ),
    .A1(\r1.regblock[29][14] ),
    .A2(\r1.regblock[30][14] ),
    .A3(\r1.regblock[31][14] ),
    .S0(net22),
    .S1(net16),
    .X(_01002_));
 sky130_fd_sc_hd__mux4_1 _13831_ (.A0(_00999_),
    .A1(_01000_),
    .A2(_01001_),
    .A3(_01002_),
    .S0(net15),
    .S1(net13),
    .X(_01003_));
 sky130_fd_sc_hd__mux4_1 _13832_ (.A0(\r1.regblock[0][13] ),
    .A1(\r1.regblock[1][13] ),
    .A2(\r1.regblock[2][13] ),
    .A3(\r1.regblock[3][13] ),
    .S0(net22),
    .S1(net16),
    .X(_00982_));
 sky130_fd_sc_hd__mux4_2 _13833_ (.A0(\r1.regblock[4][13] ),
    .A1(\r1.regblock[5][13] ),
    .A2(\r1.regblock[6][13] ),
    .A3(\r1.regblock[7][13] ),
    .S0(net24),
    .S1(net16),
    .X(_00983_));
 sky130_fd_sc_hd__mux4_1 _13834_ (.A0(\r1.regblock[8][13] ),
    .A1(\r1.regblock[9][13] ),
    .A2(\r1.regblock[10][13] ),
    .A3(\r1.regblock[11][13] ),
    .S0(net22),
    .S1(net16),
    .X(_00984_));
 sky130_fd_sc_hd__mux4_2 _13835_ (.A0(\r1.regblock[12][13] ),
    .A1(\r1.regblock[13][13] ),
    .A2(\r1.regblock[14][13] ),
    .A3(\r1.regblock[15][13] ),
    .S0(net24),
    .S1(net16),
    .X(_00985_));
 sky130_fd_sc_hd__mux4_2 _13836_ (.A0(_00982_),
    .A1(_00983_),
    .A2(_00984_),
    .A3(_00985_),
    .S0(net15),
    .S1(net13),
    .X(_00986_));
 sky130_fd_sc_hd__mux4_2 _13837_ (.A0(\r1.regblock[16][13] ),
    .A1(\r1.regblock[17][13] ),
    .A2(\r1.regblock[18][13] ),
    .A3(\r1.regblock[19][13] ),
    .S0(net22),
    .S1(net16),
    .X(_00987_));
 sky130_fd_sc_hd__mux4_2 _13838_ (.A0(\r1.regblock[20][13] ),
    .A1(\r1.regblock[21][13] ),
    .A2(\r1.regblock[22][13] ),
    .A3(\r1.regblock[23][13] ),
    .S0(net22),
    .S1(net16),
    .X(_00988_));
 sky130_fd_sc_hd__mux4_1 _13839_ (.A0(\r1.regblock[24][13] ),
    .A1(\r1.regblock[25][13] ),
    .A2(\r1.regblock[26][13] ),
    .A3(\r1.regblock[27][13] ),
    .S0(net22),
    .S1(net16),
    .X(_00989_));
 sky130_fd_sc_hd__mux4_2 _13840_ (.A0(\r1.regblock[28][13] ),
    .A1(\r1.regblock[29][13] ),
    .A2(\r1.regblock[30][13] ),
    .A3(\r1.regblock[31][13] ),
    .S0(net22),
    .S1(net16),
    .X(_00990_));
 sky130_fd_sc_hd__mux4_1 _13841_ (.A0(_00987_),
    .A1(_00988_),
    .A2(_00989_),
    .A3(_00990_),
    .S0(net15),
    .S1(net13),
    .X(_00991_));
 sky130_fd_sc_hd__mux4_2 _13842_ (.A0(\r1.regblock[0][12] ),
    .A1(\r1.regblock[1][12] ),
    .A2(\r1.regblock[2][12] ),
    .A3(\r1.regblock[3][12] ),
    .S0(net22),
    .S1(net16),
    .X(_00970_));
 sky130_fd_sc_hd__mux4_2 _13843_ (.A0(\r1.regblock[4][12] ),
    .A1(\r1.regblock[5][12] ),
    .A2(\r1.regblock[6][12] ),
    .A3(\r1.regblock[7][12] ),
    .S0(net24),
    .S1(net16),
    .X(_00971_));
 sky130_fd_sc_hd__mux4_1 _13844_ (.A0(\r1.regblock[8][12] ),
    .A1(\r1.regblock[9][12] ),
    .A2(\r1.regblock[10][12] ),
    .A3(\r1.regblock[11][12] ),
    .S0(net22),
    .S1(net16),
    .X(_00972_));
 sky130_fd_sc_hd__mux4_2 _13845_ (.A0(\r1.regblock[12][12] ),
    .A1(\r1.regblock[13][12] ),
    .A2(\r1.regblock[14][12] ),
    .A3(\r1.regblock[15][12] ),
    .S0(net24),
    .S1(net16),
    .X(_00973_));
 sky130_fd_sc_hd__mux4_2 _13846_ (.A0(_00970_),
    .A1(_00971_),
    .A2(_00972_),
    .A3(_00973_),
    .S0(net15),
    .S1(net13),
    .X(_00974_));
 sky130_fd_sc_hd__mux4_2 _13847_ (.A0(\r1.regblock[16][12] ),
    .A1(\r1.regblock[17][12] ),
    .A2(\r1.regblock[18][12] ),
    .A3(\r1.regblock[19][12] ),
    .S0(net22),
    .S1(net16),
    .X(_00975_));
 sky130_fd_sc_hd__mux4_2 _13848_ (.A0(\r1.regblock[20][12] ),
    .A1(\r1.regblock[21][12] ),
    .A2(\r1.regblock[22][12] ),
    .A3(\r1.regblock[23][12] ),
    .S0(net22),
    .S1(net16),
    .X(_00976_));
 sky130_fd_sc_hd__mux4_1 _13849_ (.A0(\r1.regblock[24][12] ),
    .A1(\r1.regblock[25][12] ),
    .A2(\r1.regblock[26][12] ),
    .A3(\r1.regblock[27][12] ),
    .S0(net22),
    .S1(net16),
    .X(_00977_));
 sky130_fd_sc_hd__mux4_1 _13850_ (.A0(\r1.regblock[28][12] ),
    .A1(\r1.regblock[29][12] ),
    .A2(\r1.regblock[30][12] ),
    .A3(\r1.regblock[31][12] ),
    .S0(net22),
    .S1(net16),
    .X(_00978_));
 sky130_fd_sc_hd__mux4_1 _13851_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00977_),
    .A3(_00978_),
    .S0(net15),
    .S1(net13),
    .X(_00979_));
 sky130_fd_sc_hd__mux4_2 _13852_ (.A0(\r1.regblock[0][11] ),
    .A1(\r1.regblock[1][11] ),
    .A2(\r1.regblock[2][11] ),
    .A3(\r1.regblock[3][11] ),
    .S0(net22),
    .S1(net16),
    .X(_00958_));
 sky130_fd_sc_hd__mux4_2 _13853_ (.A0(\r1.regblock[4][11] ),
    .A1(\r1.regblock[5][11] ),
    .A2(\r1.regblock[6][11] ),
    .A3(\r1.regblock[7][11] ),
    .S0(net24),
    .S1(net16),
    .X(_00959_));
 sky130_fd_sc_hd__mux4_1 _13854_ (.A0(\r1.regblock[8][11] ),
    .A1(\r1.regblock[9][11] ),
    .A2(\r1.regblock[10][11] ),
    .A3(\r1.regblock[11][11] ),
    .S0(net24),
    .S1(net16),
    .X(_00960_));
 sky130_fd_sc_hd__mux4_1 _13855_ (.A0(\r1.regblock[12][11] ),
    .A1(\r1.regblock[13][11] ),
    .A2(\r1.regblock[14][11] ),
    .A3(\r1.regblock[15][11] ),
    .S0(net24),
    .S1(net16),
    .X(_00961_));
 sky130_fd_sc_hd__mux4_2 _13856_ (.A0(_00958_),
    .A1(_00959_),
    .A2(_00960_),
    .A3(_00961_),
    .S0(net15),
    .S1(net13),
    .X(_00962_));
 sky130_fd_sc_hd__mux4_2 _13857_ (.A0(\r1.regblock[16][11] ),
    .A1(\r1.regblock[17][11] ),
    .A2(\r1.regblock[18][11] ),
    .A3(\r1.regblock[19][11] ),
    .S0(net22),
    .S1(net16),
    .X(_00963_));
 sky130_fd_sc_hd__mux4_2 _13858_ (.A0(\r1.regblock[20][11] ),
    .A1(\r1.regblock[21][11] ),
    .A2(\r1.regblock[22][11] ),
    .A3(\r1.regblock[23][11] ),
    .S0(net22),
    .S1(net16),
    .X(_00964_));
 sky130_fd_sc_hd__mux4_2 _13859_ (.A0(\r1.regblock[24][11] ),
    .A1(\r1.regblock[25][11] ),
    .A2(\r1.regblock[26][11] ),
    .A3(\r1.regblock[27][11] ),
    .S0(net22),
    .S1(net16),
    .X(_00965_));
 sky130_fd_sc_hd__mux4_2 _13860_ (.A0(\r1.regblock[28][11] ),
    .A1(\r1.regblock[29][11] ),
    .A2(\r1.regblock[30][11] ),
    .A3(\r1.regblock[31][11] ),
    .S0(net22),
    .S1(net16),
    .X(_00966_));
 sky130_fd_sc_hd__mux4_1 _13861_ (.A0(_00963_),
    .A1(_00964_),
    .A2(_00965_),
    .A3(_00966_),
    .S0(net15),
    .S1(net13),
    .X(_00967_));
 sky130_fd_sc_hd__mux4_1 _13862_ (.A0(\r1.regblock[0][10] ),
    .A1(\r1.regblock[1][10] ),
    .A2(\r1.regblock[2][10] ),
    .A3(\r1.regblock[3][10] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00946_));
 sky130_fd_sc_hd__mux4_2 _13863_ (.A0(\r1.regblock[4][10] ),
    .A1(\r1.regblock[5][10] ),
    .A2(\r1.regblock[6][10] ),
    .A3(\r1.regblock[7][10] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00947_));
 sky130_fd_sc_hd__mux4_1 _13864_ (.A0(\r1.regblock[8][10] ),
    .A1(\r1.regblock[9][10] ),
    .A2(\r1.regblock[10][10] ),
    .A3(\r1.regblock[11][10] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00948_));
 sky130_fd_sc_hd__mux4_1 _13865_ (.A0(\r1.regblock[12][10] ),
    .A1(\r1.regblock[13][10] ),
    .A2(\r1.regblock[14][10] ),
    .A3(\r1.regblock[15][10] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00949_));
 sky130_fd_sc_hd__mux4_2 _13866_ (.A0(_00946_),
    .A1(_00947_),
    .A2(_00948_),
    .A3(_00949_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00950_));
 sky130_fd_sc_hd__mux4_2 _13867_ (.A0(\r1.regblock[16][10] ),
    .A1(\r1.regblock[17][10] ),
    .A2(\r1.regblock[18][10] ),
    .A3(\r1.regblock[19][10] ),
    .S0(net30),
    .S1(net21),
    .X(_00951_));
 sky130_fd_sc_hd__mux4_1 _13868_ (.A0(\r1.regblock[20][10] ),
    .A1(\r1.regblock[21][10] ),
    .A2(\r1.regblock[22][10] ),
    .A3(\r1.regblock[23][10] ),
    .S0(net30),
    .S1(net21),
    .X(_00952_));
 sky130_fd_sc_hd__mux4_1 _13869_ (.A0(\r1.regblock[24][10] ),
    .A1(\r1.regblock[25][10] ),
    .A2(\r1.regblock[26][10] ),
    .A3(\r1.regblock[27][10] ),
    .S0(net30),
    .S1(net21),
    .X(_00953_));
 sky130_fd_sc_hd__mux4_2 _13870_ (.A0(\r1.regblock[28][10] ),
    .A1(\r1.regblock[29][10] ),
    .A2(\r1.regblock[30][10] ),
    .A3(\r1.regblock[31][10] ),
    .S0(net30),
    .S1(net21),
    .X(_00954_));
 sky130_fd_sc_hd__mux4_2 _13871_ (.A0(_00951_),
    .A1(_00952_),
    .A2(_00953_),
    .A3(_00954_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00955_));
 sky130_fd_sc_hd__mux4_1 _13872_ (.A0(\r1.regblock[0][9] ),
    .A1(\r1.regblock[1][9] ),
    .A2(\r1.regblock[2][9] ),
    .A3(\r1.regblock[3][9] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00934_));
 sky130_fd_sc_hd__mux4_2 _13873_ (.A0(\r1.regblock[4][9] ),
    .A1(\r1.regblock[5][9] ),
    .A2(\r1.regblock[6][9] ),
    .A3(\r1.regblock[7][9] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00935_));
 sky130_fd_sc_hd__mux4_2 _13874_ (.A0(\r1.regblock[8][9] ),
    .A1(\r1.regblock[9][9] ),
    .A2(\r1.regblock[10][9] ),
    .A3(\r1.regblock[11][9] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00936_));
 sky130_fd_sc_hd__mux4_1 _13875_ (.A0(\r1.regblock[12][9] ),
    .A1(\r1.regblock[13][9] ),
    .A2(\r1.regblock[14][9] ),
    .A3(\r1.regblock[15][9] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00937_));
 sky130_fd_sc_hd__mux4_2 _13876_ (.A0(_00934_),
    .A1(_00935_),
    .A2(_00936_),
    .A3(_00937_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00938_));
 sky130_fd_sc_hd__mux4_1 _13877_ (.A0(\r1.regblock[16][9] ),
    .A1(\r1.regblock[17][9] ),
    .A2(\r1.regblock[18][9] ),
    .A3(\r1.regblock[19][9] ),
    .S0(net30),
    .S1(net21),
    .X(_00939_));
 sky130_fd_sc_hd__mux4_2 _13878_ (.A0(\r1.regblock[20][9] ),
    .A1(\r1.regblock[21][9] ),
    .A2(\r1.regblock[22][9] ),
    .A3(\r1.regblock[23][9] ),
    .S0(net30),
    .S1(net21),
    .X(_00940_));
 sky130_fd_sc_hd__mux4_1 _13879_ (.A0(\r1.regblock[24][9] ),
    .A1(\r1.regblock[25][9] ),
    .A2(\r1.regblock[26][9] ),
    .A3(\r1.regblock[27][9] ),
    .S0(net30),
    .S1(net21),
    .X(_00941_));
 sky130_fd_sc_hd__mux4_2 _13880_ (.A0(\r1.regblock[28][9] ),
    .A1(\r1.regblock[29][9] ),
    .A2(\r1.regblock[30][9] ),
    .A3(\r1.regblock[31][9] ),
    .S0(net30),
    .S1(net21),
    .X(_00942_));
 sky130_fd_sc_hd__mux4_2 _13881_ (.A0(_00939_),
    .A1(_00940_),
    .A2(_00941_),
    .A3(_00942_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00943_));
 sky130_fd_sc_hd__mux4_1 _13882_ (.A0(\r1.regblock[0][8] ),
    .A1(\r1.regblock[1][8] ),
    .A2(\r1.regblock[2][8] ),
    .A3(\r1.regblock[3][8] ),
    .S0(net30),
    .S1(net21),
    .X(_00922_));
 sky130_fd_sc_hd__mux4_2 _13883_ (.A0(\r1.regblock[4][8] ),
    .A1(\r1.regblock[5][8] ),
    .A2(\r1.regblock[6][8] ),
    .A3(\r1.regblock[7][8] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00923_));
 sky130_fd_sc_hd__mux4_2 _13884_ (.A0(\r1.regblock[8][8] ),
    .A1(\r1.regblock[9][8] ),
    .A2(\r1.regblock[10][8] ),
    .A3(\r1.regblock[11][8] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00924_));
 sky130_fd_sc_hd__mux4_2 _13885_ (.A0(\r1.regblock[12][8] ),
    .A1(\r1.regblock[13][8] ),
    .A2(\r1.regblock[14][8] ),
    .A3(\r1.regblock[15][8] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00925_));
 sky130_fd_sc_hd__mux4_2 _13886_ (.A0(_00922_),
    .A1(_00923_),
    .A2(_00924_),
    .A3(_00925_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00926_));
 sky130_fd_sc_hd__mux4_1 _13887_ (.A0(\r1.regblock[16][8] ),
    .A1(\r1.regblock[17][8] ),
    .A2(\r1.regblock[18][8] ),
    .A3(\r1.regblock[19][8] ),
    .S0(net30),
    .S1(net21),
    .X(_00927_));
 sky130_fd_sc_hd__mux4_2 _13888_ (.A0(\r1.regblock[20][8] ),
    .A1(\r1.regblock[21][8] ),
    .A2(\r1.regblock[22][8] ),
    .A3(\r1.regblock[23][8] ),
    .S0(net30),
    .S1(net21),
    .X(_00928_));
 sky130_fd_sc_hd__mux4_1 _13889_ (.A0(\r1.regblock[24][8] ),
    .A1(\r1.regblock[25][8] ),
    .A2(\r1.regblock[26][8] ),
    .A3(\r1.regblock[27][8] ),
    .S0(net30),
    .S1(net21),
    .X(_00929_));
 sky130_fd_sc_hd__mux4_2 _13890_ (.A0(\r1.regblock[28][8] ),
    .A1(\r1.regblock[29][8] ),
    .A2(\r1.regblock[30][8] ),
    .A3(\r1.regblock[31][8] ),
    .S0(net30),
    .S1(net21),
    .X(_00930_));
 sky130_fd_sc_hd__mux4_2 _13891_ (.A0(_00927_),
    .A1(_00928_),
    .A2(_00929_),
    .A3(_00930_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00931_));
 sky130_fd_sc_hd__mux4_2 _13892_ (.A0(\r1.regblock[0][7] ),
    .A1(\r1.regblock[1][7] ),
    .A2(\r1.regblock[2][7] ),
    .A3(\r1.regblock[3][7] ),
    .S0(net30),
    .S1(net21),
    .X(_00910_));
 sky130_fd_sc_hd__mux4_2 _13893_ (.A0(\r1.regblock[4][7] ),
    .A1(\r1.regblock[5][7] ),
    .A2(\r1.regblock[6][7] ),
    .A3(\r1.regblock[7][7] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00911_));
 sky130_fd_sc_hd__mux4_1 _13894_ (.A0(\r1.regblock[8][7] ),
    .A1(\r1.regblock[9][7] ),
    .A2(\r1.regblock[10][7] ),
    .A3(\r1.regblock[11][7] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00912_));
 sky130_fd_sc_hd__mux4_1 _13895_ (.A0(\r1.regblock[12][7] ),
    .A1(\r1.regblock[13][7] ),
    .A2(\r1.regblock[14][7] ),
    .A3(\r1.regblock[15][7] ),
    .S0(\c1.instruction1[15] ),
    .S1(\c1.instruction1[16] ),
    .X(_00913_));
 sky130_fd_sc_hd__mux4_2 _13896_ (.A0(_00910_),
    .A1(_00911_),
    .A2(_00912_),
    .A3(_00913_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00914_));
 sky130_fd_sc_hd__mux4_1 _13897_ (.A0(\r1.regblock[16][7] ),
    .A1(\r1.regblock[17][7] ),
    .A2(\r1.regblock[18][7] ),
    .A3(\r1.regblock[19][7] ),
    .S0(net29),
    .S1(net21),
    .X(_00915_));
 sky130_fd_sc_hd__mux4_2 _13898_ (.A0(\r1.regblock[20][7] ),
    .A1(\r1.regblock[21][7] ),
    .A2(\r1.regblock[22][7] ),
    .A3(\r1.regblock[23][7] ),
    .S0(net30),
    .S1(net21),
    .X(_00916_));
 sky130_fd_sc_hd__mux4_2 _13899_ (.A0(\r1.regblock[24][7] ),
    .A1(\r1.regblock[25][7] ),
    .A2(\r1.regblock[26][7] ),
    .A3(\r1.regblock[27][7] ),
    .S0(net30),
    .S1(net21),
    .X(_00917_));
 sky130_fd_sc_hd__mux4_2 _13900_ (.A0(\r1.regblock[28][7] ),
    .A1(\r1.regblock[29][7] ),
    .A2(\r1.regblock[30][7] ),
    .A3(\r1.regblock[31][7] ),
    .S0(net30),
    .S1(net21),
    .X(_00918_));
 sky130_fd_sc_hd__mux4_1 _13901_ (.A0(_00915_),
    .A1(_00916_),
    .A2(_00917_),
    .A3(_00918_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00919_));
 sky130_fd_sc_hd__mux4_1 _13902_ (.A0(\r1.regblock[0][6] ),
    .A1(\r1.regblock[1][6] ),
    .A2(\r1.regblock[2][6] ),
    .A3(\r1.regblock[3][6] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00898_));
 sky130_fd_sc_hd__mux4_2 _13903_ (.A0(\r1.regblock[4][6] ),
    .A1(\r1.regblock[5][6] ),
    .A2(\r1.regblock[6][6] ),
    .A3(\r1.regblock[7][6] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00899_));
 sky130_fd_sc_hd__mux4_2 _13904_ (.A0(\r1.regblock[8][6] ),
    .A1(\r1.regblock[9][6] ),
    .A2(\r1.regblock[10][6] ),
    .A3(\r1.regblock[11][6] ),
    .S0(net30),
    .S1(net21),
    .X(_00900_));
 sky130_fd_sc_hd__mux4_1 _13905_ (.A0(\r1.regblock[12][6] ),
    .A1(\r1.regblock[13][6] ),
    .A2(\r1.regblock[14][6] ),
    .A3(\r1.regblock[15][6] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00901_));
 sky130_fd_sc_hd__mux4_2 _13906_ (.A0(_00898_),
    .A1(_00899_),
    .A2(_00900_),
    .A3(_00901_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00902_));
 sky130_fd_sc_hd__mux4_1 _13907_ (.A0(\r1.regblock[16][6] ),
    .A1(\r1.regblock[17][6] ),
    .A2(\r1.regblock[18][6] ),
    .A3(\r1.regblock[19][6] ),
    .S0(net29),
    .S1(net21),
    .X(_00903_));
 sky130_fd_sc_hd__mux4_2 _13908_ (.A0(\r1.regblock[20][6] ),
    .A1(\r1.regblock[21][6] ),
    .A2(\r1.regblock[22][6] ),
    .A3(\r1.regblock[23][6] ),
    .S0(net24),
    .S1(net17),
    .X(_00904_));
 sky130_fd_sc_hd__mux4_2 _13909_ (.A0(\r1.regblock[24][6] ),
    .A1(\r1.regblock[25][6] ),
    .A2(\r1.regblock[26][6] ),
    .A3(\r1.regblock[27][6] ),
    .S0(net30),
    .S1(net21),
    .X(_00905_));
 sky130_fd_sc_hd__mux4_1 _13910_ (.A0(\r1.regblock[28][6] ),
    .A1(\r1.regblock[29][6] ),
    .A2(\r1.regblock[30][6] ),
    .A3(\r1.regblock[31][6] ),
    .S0(net29),
    .S1(net21),
    .X(_00906_));
 sky130_fd_sc_hd__mux4_1 _13911_ (.A0(_00903_),
    .A1(_00904_),
    .A2(_00905_),
    .A3(_00906_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00907_));
 sky130_fd_sc_hd__mux4_2 _13912_ (.A0(\r1.regblock[0][5] ),
    .A1(\r1.regblock[1][5] ),
    .A2(\r1.regblock[2][5] ),
    .A3(\r1.regblock[3][5] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00886_));
 sky130_fd_sc_hd__mux4_2 _13913_ (.A0(\r1.regblock[4][5] ),
    .A1(\r1.regblock[5][5] ),
    .A2(\r1.regblock[6][5] ),
    .A3(\r1.regblock[7][5] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00887_));
 sky130_fd_sc_hd__mux4_1 _13914_ (.A0(\r1.regblock[8][5] ),
    .A1(\r1.regblock[9][5] ),
    .A2(\r1.regblock[10][5] ),
    .A3(\r1.regblock[11][5] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00888_));
 sky130_fd_sc_hd__mux4_1 _13915_ (.A0(\r1.regblock[12][5] ),
    .A1(\r1.regblock[13][5] ),
    .A2(\r1.regblock[14][5] ),
    .A3(\r1.regblock[15][5] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00889_));
 sky130_fd_sc_hd__mux4_2 _13916_ (.A0(_00886_),
    .A1(_00887_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00890_));
 sky130_fd_sc_hd__mux4_1 _13917_ (.A0(\r1.regblock[16][5] ),
    .A1(\r1.regblock[17][5] ),
    .A2(\r1.regblock[18][5] ),
    .A3(\r1.regblock[19][5] ),
    .S0(net29),
    .S1(net21),
    .X(_00891_));
 sky130_fd_sc_hd__mux4_2 _13918_ (.A0(\r1.regblock[20][5] ),
    .A1(\r1.regblock[21][5] ),
    .A2(\r1.regblock[22][5] ),
    .A3(\r1.regblock[23][5] ),
    .S0(net24),
    .S1(net17),
    .X(_00892_));
 sky130_fd_sc_hd__mux4_2 _13919_ (.A0(\r1.regblock[24][5] ),
    .A1(\r1.regblock[25][5] ),
    .A2(\r1.regblock[26][5] ),
    .A3(\r1.regblock[27][5] ),
    .S0(net30),
    .S1(net21),
    .X(_00893_));
 sky130_fd_sc_hd__mux4_2 _13920_ (.A0(\r1.regblock[28][5] ),
    .A1(\r1.regblock[29][5] ),
    .A2(\r1.regblock[30][5] ),
    .A3(\r1.regblock[31][5] ),
    .S0(net29),
    .S1(net21),
    .X(_00894_));
 sky130_fd_sc_hd__mux4_1 _13921_ (.A0(_00891_),
    .A1(_00892_),
    .A2(_00893_),
    .A3(_00894_),
    .S0(\c1.instruction1[17] ),
    .S1(net12),
    .X(_00895_));
 sky130_fd_sc_hd__mux4_2 _13922_ (.A0(\r1.regblock[0][4] ),
    .A1(\r1.regblock[1][4] ),
    .A2(\r1.regblock[2][4] ),
    .A3(\r1.regblock[3][4] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00874_));
 sky130_fd_sc_hd__mux4_2 _13923_ (.A0(\r1.regblock[4][4] ),
    .A1(\r1.regblock[5][4] ),
    .A2(\r1.regblock[6][4] ),
    .A3(\r1.regblock[7][4] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00875_));
 sky130_fd_sc_hd__mux4_1 _13924_ (.A0(\r1.regblock[8][4] ),
    .A1(\r1.regblock[9][4] ),
    .A2(\r1.regblock[10][4] ),
    .A3(\r1.regblock[11][4] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00876_));
 sky130_fd_sc_hd__mux4_1 _13925_ (.A0(\r1.regblock[12][4] ),
    .A1(\r1.regblock[13][4] ),
    .A2(\r1.regblock[14][4] ),
    .A3(\r1.regblock[15][4] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00877_));
 sky130_fd_sc_hd__mux4_2 _13926_ (.A0(_00874_),
    .A1(_00875_),
    .A2(_00876_),
    .A3(_00877_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00878_));
 sky130_fd_sc_hd__mux4_1 _13927_ (.A0(\r1.regblock[16][4] ),
    .A1(\r1.regblock[17][4] ),
    .A2(\r1.regblock[18][4] ),
    .A3(\r1.regblock[19][4] ),
    .S0(net29),
    .S1(net21),
    .X(_00879_));
 sky130_fd_sc_hd__mux4_2 _13928_ (.A0(\r1.regblock[20][4] ),
    .A1(\r1.regblock[21][4] ),
    .A2(\r1.regblock[22][4] ),
    .A3(\r1.regblock[23][4] ),
    .S0(net29),
    .S1(net21),
    .X(_00880_));
 sky130_fd_sc_hd__mux4_1 _13929_ (.A0(\r1.regblock[24][4] ),
    .A1(\r1.regblock[25][4] ),
    .A2(\r1.regblock[26][4] ),
    .A3(\r1.regblock[27][4] ),
    .S0(net29),
    .S1(net21),
    .X(_00881_));
 sky130_fd_sc_hd__mux4_2 _13930_ (.A0(\r1.regblock[28][4] ),
    .A1(\r1.regblock[29][4] ),
    .A2(\r1.regblock[30][4] ),
    .A3(\r1.regblock[31][4] ),
    .S0(net29),
    .S1(net21),
    .X(_00882_));
 sky130_fd_sc_hd__mux4_1 _13931_ (.A0(_00879_),
    .A1(_00880_),
    .A2(_00881_),
    .A3(_00882_),
    .S0(\c1.instruction1[17] ),
    .S1(net12),
    .X(_00883_));
 sky130_fd_sc_hd__mux4_2 _13932_ (.A0(\r1.regblock[0][3] ),
    .A1(\r1.regblock[1][3] ),
    .A2(\r1.regblock[2][3] ),
    .A3(\r1.regblock[3][3] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00862_));
 sky130_fd_sc_hd__mux4_2 _13933_ (.A0(\r1.regblock[4][3] ),
    .A1(\r1.regblock[5][3] ),
    .A2(\r1.regblock[6][3] ),
    .A3(\r1.regblock[7][3] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00863_));
 sky130_fd_sc_hd__mux4_1 _13934_ (.A0(\r1.regblock[8][3] ),
    .A1(\r1.regblock[9][3] ),
    .A2(\r1.regblock[10][3] ),
    .A3(\r1.regblock[11][3] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00864_));
 sky130_fd_sc_hd__mux4_1 _13935_ (.A0(\r1.regblock[12][3] ),
    .A1(\r1.regblock[13][3] ),
    .A2(\r1.regblock[14][3] ),
    .A3(\r1.regblock[15][3] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00865_));
 sky130_fd_sc_hd__mux4_2 _13936_ (.A0(_00862_),
    .A1(_00863_),
    .A2(_00864_),
    .A3(_00865_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00866_));
 sky130_fd_sc_hd__mux4_1 _13937_ (.A0(\r1.regblock[16][3] ),
    .A1(\r1.regblock[17][3] ),
    .A2(\r1.regblock[18][3] ),
    .A3(\r1.regblock[19][3] ),
    .S0(net28),
    .S1(net21),
    .X(_00867_));
 sky130_fd_sc_hd__mux4_2 _13938_ (.A0(\r1.regblock[20][3] ),
    .A1(\r1.regblock[21][3] ),
    .A2(\r1.regblock[22][3] ),
    .A3(\r1.regblock[23][3] ),
    .S0(net29),
    .S1(net21),
    .X(_00868_));
 sky130_fd_sc_hd__mux4_1 _13939_ (.A0(\r1.regblock[24][3] ),
    .A1(\r1.regblock[25][3] ),
    .A2(\r1.regblock[26][3] ),
    .A3(\r1.regblock[27][3] ),
    .S0(net29),
    .S1(net21),
    .X(_00869_));
 sky130_fd_sc_hd__mux4_2 _13940_ (.A0(\r1.regblock[28][3] ),
    .A1(\r1.regblock[29][3] ),
    .A2(\r1.regblock[30][3] ),
    .A3(\r1.regblock[31][3] ),
    .S0(net29),
    .S1(net21),
    .X(_00870_));
 sky130_fd_sc_hd__mux4_1 _13941_ (.A0(_00867_),
    .A1(_00868_),
    .A2(_00869_),
    .A3(_00870_),
    .S0(net14),
    .S1(net12),
    .X(_00871_));
 sky130_fd_sc_hd__mux4_2 _13942_ (.A0(\r1.regblock[0][2] ),
    .A1(\r1.regblock[1][2] ),
    .A2(\r1.regblock[2][2] ),
    .A3(\r1.regblock[3][2] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00850_));
 sky130_fd_sc_hd__mux4_2 _13943_ (.A0(\r1.regblock[4][2] ),
    .A1(\r1.regblock[5][2] ),
    .A2(\r1.regblock[6][2] ),
    .A3(\r1.regblock[7][2] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00851_));
 sky130_fd_sc_hd__mux4_1 _13944_ (.A0(\r1.regblock[8][2] ),
    .A1(\r1.regblock[9][2] ),
    .A2(\r1.regblock[10][2] ),
    .A3(\r1.regblock[11][2] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00852_));
 sky130_fd_sc_hd__mux4_2 _13945_ (.A0(\r1.regblock[12][2] ),
    .A1(\r1.regblock[13][2] ),
    .A2(\r1.regblock[14][2] ),
    .A3(\r1.regblock[15][2] ),
    .S0(net31),
    .S1(\c1.instruction1[16] ),
    .X(_00853_));
 sky130_fd_sc_hd__mux4_2 _13946_ (.A0(_00850_),
    .A1(_00851_),
    .A2(_00852_),
    .A3(_00853_),
    .S0(\c1.instruction1[17] ),
    .S1(net13),
    .X(_00854_));
 sky130_fd_sc_hd__mux4_1 _13947_ (.A0(\r1.regblock[16][2] ),
    .A1(\r1.regblock[17][2] ),
    .A2(\r1.regblock[18][2] ),
    .A3(\r1.regblock[19][2] ),
    .S0(net28),
    .S1(net20),
    .X(_00855_));
 sky130_fd_sc_hd__mux4_2 _13948_ (.A0(\r1.regblock[20][2] ),
    .A1(\r1.regblock[21][2] ),
    .A2(\r1.regblock[22][2] ),
    .A3(\r1.regblock[23][2] ),
    .S0(net29),
    .S1(net21),
    .X(_00856_));
 sky130_fd_sc_hd__mux4_1 _13949_ (.A0(\r1.regblock[24][2] ),
    .A1(\r1.regblock[25][2] ),
    .A2(\r1.regblock[26][2] ),
    .A3(\r1.regblock[27][2] ),
    .S0(net29),
    .S1(net21),
    .X(_00857_));
 sky130_fd_sc_hd__mux4_2 _13950_ (.A0(\r1.regblock[28][2] ),
    .A1(\r1.regblock[29][2] ),
    .A2(\r1.regblock[30][2] ),
    .A3(\r1.regblock[31][2] ),
    .S0(net29),
    .S1(net21),
    .X(_00858_));
 sky130_fd_sc_hd__mux4_1 _13951_ (.A0(_00855_),
    .A1(_00856_),
    .A2(_00857_),
    .A3(_00858_),
    .S0(net14),
    .S1(net12),
    .X(_00859_));
 sky130_fd_sc_hd__mux4_2 _13952_ (.A0(\r1.regblock[0][1] ),
    .A1(\r1.regblock[1][1] ),
    .A2(\r1.regblock[2][1] ),
    .A3(\r1.regblock[3][1] ),
    .S0(net28),
    .S1(net20),
    .X(_00838_));
 sky130_fd_sc_hd__mux4_2 _13953_ (.A0(\r1.regblock[4][1] ),
    .A1(\r1.regblock[5][1] ),
    .A2(\r1.regblock[6][1] ),
    .A3(\r1.regblock[7][1] ),
    .S0(net25),
    .S1(net18),
    .X(_00839_));
 sky130_fd_sc_hd__mux4_1 _13954_ (.A0(\r1.regblock[8][1] ),
    .A1(\r1.regblock[9][1] ),
    .A2(\r1.regblock[10][1] ),
    .A3(\r1.regblock[11][1] ),
    .S0(net28),
    .S1(net20),
    .X(_00840_));
 sky130_fd_sc_hd__mux4_1 _13955_ (.A0(\r1.regblock[12][1] ),
    .A1(\r1.regblock[13][1] ),
    .A2(\r1.regblock[14][1] ),
    .A3(\r1.regblock[15][1] ),
    .S0(net28),
    .S1(net20),
    .X(_00841_));
 sky130_fd_sc_hd__mux4_2 _13956_ (.A0(_00838_),
    .A1(_00839_),
    .A2(_00840_),
    .A3(_00841_),
    .S0(net14),
    .S1(net12),
    .X(_00842_));
 sky130_fd_sc_hd__mux4_2 _13957_ (.A0(\r1.regblock[16][1] ),
    .A1(\r1.regblock[17][1] ),
    .A2(\r1.regblock[18][1] ),
    .A3(\r1.regblock[19][1] ),
    .S0(net28),
    .S1(net20),
    .X(_00843_));
 sky130_fd_sc_hd__mux4_2 _13958_ (.A0(\r1.regblock[20][1] ),
    .A1(\r1.regblock[21][1] ),
    .A2(\r1.regblock[22][1] ),
    .A3(\r1.regblock[23][1] ),
    .S0(net28),
    .S1(net20),
    .X(_00844_));
 sky130_fd_sc_hd__mux4_1 _13959_ (.A0(\r1.regblock[24][1] ),
    .A1(\r1.regblock[25][1] ),
    .A2(\r1.regblock[26][1] ),
    .A3(\r1.regblock[27][1] ),
    .S0(net28),
    .S1(net20),
    .X(_00845_));
 sky130_fd_sc_hd__mux4_2 _13960_ (.A0(\r1.regblock[28][1] ),
    .A1(\r1.regblock[29][1] ),
    .A2(\r1.regblock[30][1] ),
    .A3(\r1.regblock[31][1] ),
    .S0(net28),
    .S1(net20),
    .X(_00846_));
 sky130_fd_sc_hd__mux4_1 _13961_ (.A0(_00843_),
    .A1(_00844_),
    .A2(_00845_),
    .A3(_00846_),
    .S0(net15),
    .S1(\c1.instruction1[18] ),
    .X(_00847_));
 sky130_fd_sc_hd__mux4_2 _13962_ (.A0(\r1.regblock[0][0] ),
    .A1(\r1.regblock[1][0] ),
    .A2(\r1.regblock[2][0] ),
    .A3(\r1.regblock[3][0] ),
    .S0(net28),
    .S1(net20),
    .X(_00826_));
 sky130_fd_sc_hd__mux4_2 _13963_ (.A0(\r1.regblock[4][0] ),
    .A1(\r1.regblock[5][0] ),
    .A2(\r1.regblock[6][0] ),
    .A3(\r1.regblock[7][0] ),
    .S0(net25),
    .S1(net18),
    .X(_00827_));
 sky130_fd_sc_hd__mux4_1 _13964_ (.A0(\r1.regblock[8][0] ),
    .A1(\r1.regblock[9][0] ),
    .A2(\r1.regblock[10][0] ),
    .A3(\r1.regblock[11][0] ),
    .S0(net28),
    .S1(net20),
    .X(_00828_));
 sky130_fd_sc_hd__mux4_1 _13965_ (.A0(\r1.regblock[12][0] ),
    .A1(\r1.regblock[13][0] ),
    .A2(\r1.regblock[14][0] ),
    .A3(\r1.regblock[15][0] ),
    .S0(net28),
    .S1(net20),
    .X(_00829_));
 sky130_fd_sc_hd__mux4_2 _13966_ (.A0(_00826_),
    .A1(_00827_),
    .A2(_00828_),
    .A3(_00829_),
    .S0(net14),
    .S1(net12),
    .X(_00830_));
 sky130_fd_sc_hd__mux4_1 _13967_ (.A0(\r1.regblock[16][0] ),
    .A1(\r1.regblock[17][0] ),
    .A2(\r1.regblock[18][0] ),
    .A3(\r1.regblock[19][0] ),
    .S0(net28),
    .S1(net20),
    .X(_00831_));
 sky130_fd_sc_hd__mux4_1 _13968_ (.A0(\r1.regblock[20][0] ),
    .A1(\r1.regblock[21][0] ),
    .A2(\r1.regblock[22][0] ),
    .A3(\r1.regblock[23][0] ),
    .S0(net28),
    .S1(net20),
    .X(_00832_));
 sky130_fd_sc_hd__mux4_1 _13969_ (.A0(\r1.regblock[24][0] ),
    .A1(\r1.regblock[25][0] ),
    .A2(\r1.regblock[26][0] ),
    .A3(\r1.regblock[27][0] ),
    .S0(net28),
    .S1(net20),
    .X(_00833_));
 sky130_fd_sc_hd__mux4_2 _13970_ (.A0(\r1.regblock[28][0] ),
    .A1(\r1.regblock[29][0] ),
    .A2(\r1.regblock[30][0] ),
    .A3(\r1.regblock[31][0] ),
    .S0(net28),
    .S1(net20),
    .X(_00834_));
 sky130_fd_sc_hd__mux4_1 _13971_ (.A0(_00831_),
    .A1(_00832_),
    .A2(_00833_),
    .A3(_00834_),
    .S0(net15),
    .S1(\c1.instruction1[18] ),
    .X(_00835_));
 sky130_fd_sc_hd__mux4_1 _13972_ (.A0(\r1.regblock[0][31] ),
    .A1(\r1.regblock[1][31] ),
    .A2(\r1.regblock[2][31] ),
    .A3(\r1.regblock[3][31] ),
    .S0(net51),
    .S1(net37),
    .X(_00813_));
 sky130_fd_sc_hd__mux4_2 _13973_ (.A0(\r1.regblock[4][31] ),
    .A1(\r1.regblock[5][31] ),
    .A2(\r1.regblock[6][31] ),
    .A3(\r1.regblock[7][31] ),
    .S0(net43),
    .S1(net38),
    .X(_00814_));
 sky130_fd_sc_hd__mux4_2 _13974_ (.A0(\r1.regblock[8][31] ),
    .A1(\r1.regblock[9][31] ),
    .A2(\r1.regblock[10][31] ),
    .A3(\r1.regblock[11][31] ),
    .S0(net51),
    .S1(net37),
    .X(_00815_));
 sky130_fd_sc_hd__mux4_1 _13975_ (.A0(\r1.regblock[12][31] ),
    .A1(\r1.regblock[13][31] ),
    .A2(\r1.regblock[14][31] ),
    .A3(\r1.regblock[15][31] ),
    .S0(net51),
    .S1(net37),
    .X(_00816_));
 sky130_fd_sc_hd__mux4_2 _13976_ (.A0(_00813_),
    .A1(_00814_),
    .A2(_00815_),
    .A3(_00816_),
    .S0(net34),
    .S1(net32),
    .X(_00817_));
 sky130_fd_sc_hd__mux4_2 _13977_ (.A0(\r1.regblock[16][31] ),
    .A1(\r1.regblock[17][31] ),
    .A2(\r1.regblock[18][31] ),
    .A3(\r1.regblock[19][31] ),
    .S0(net50),
    .S1(net37),
    .X(_00818_));
 sky130_fd_sc_hd__mux4_1 _13978_ (.A0(\r1.regblock[20][31] ),
    .A1(\r1.regblock[21][31] ),
    .A2(\r1.regblock[22][31] ),
    .A3(\r1.regblock[23][31] ),
    .S0(net50),
    .S1(net37),
    .X(_00819_));
 sky130_fd_sc_hd__mux4_1 _13979_ (.A0(\r1.regblock[24][31] ),
    .A1(\r1.regblock[25][31] ),
    .A2(\r1.regblock[26][31] ),
    .A3(\r1.regblock[27][31] ),
    .S0(net50),
    .S1(net40),
    .X(_00820_));
 sky130_fd_sc_hd__mux4_2 _13980_ (.A0(\r1.regblock[28][31] ),
    .A1(\r1.regblock[29][31] ),
    .A2(\r1.regblock[30][31] ),
    .A3(\r1.regblock[31][31] ),
    .S0(net51),
    .S1(net37),
    .X(_00821_));
 sky130_fd_sc_hd__mux4_1 _13981_ (.A0(_00818_),
    .A1(_00819_),
    .A2(_00820_),
    .A3(_00821_),
    .S0(\c1.instruction1[22] ),
    .S1(\c1.instruction1[23] ),
    .X(_00822_));
 sky130_fd_sc_hd__mux4_1 _13982_ (.A0(\r1.regblock[0][30] ),
    .A1(\r1.regblock[1][30] ),
    .A2(\r1.regblock[2][30] ),
    .A3(\r1.regblock[3][30] ),
    .S0(net51),
    .S1(net37),
    .X(_00800_));
 sky130_fd_sc_hd__mux4_2 _13983_ (.A0(\r1.regblock[4][30] ),
    .A1(\r1.regblock[5][30] ),
    .A2(\r1.regblock[6][30] ),
    .A3(\r1.regblock[7][30] ),
    .S0(net51),
    .S1(net37),
    .X(_00801_));
 sky130_fd_sc_hd__mux4_2 _13984_ (.A0(\r1.regblock[8][30] ),
    .A1(\r1.regblock[9][30] ),
    .A2(\r1.regblock[10][30] ),
    .A3(\r1.regblock[11][30] ),
    .S0(net51),
    .S1(net37),
    .X(_00802_));
 sky130_fd_sc_hd__mux4_1 _13985_ (.A0(\r1.regblock[12][30] ),
    .A1(\r1.regblock[13][30] ),
    .A2(\r1.regblock[14][30] ),
    .A3(\r1.regblock[15][30] ),
    .S0(net51),
    .S1(net37),
    .X(_00803_));
 sky130_fd_sc_hd__mux4_2 _13986_ (.A0(_00800_),
    .A1(_00801_),
    .A2(_00802_),
    .A3(_00803_),
    .S0(net34),
    .S1(net32),
    .X(_00804_));
 sky130_fd_sc_hd__mux4_1 _13987_ (.A0(\r1.regblock[16][30] ),
    .A1(\r1.regblock[17][30] ),
    .A2(\r1.regblock[18][30] ),
    .A3(\r1.regblock[19][30] ),
    .S0(net51),
    .S1(net37),
    .X(_00805_));
 sky130_fd_sc_hd__mux4_1 _13988_ (.A0(\r1.regblock[20][30] ),
    .A1(\r1.regblock[21][30] ),
    .A2(\r1.regblock[22][30] ),
    .A3(\r1.regblock[23][30] ),
    .S0(net51),
    .S1(net37),
    .X(_00806_));
 sky130_fd_sc_hd__mux4_2 _13989_ (.A0(\r1.regblock[24][30] ),
    .A1(\r1.regblock[25][30] ),
    .A2(\r1.regblock[26][30] ),
    .A3(\r1.regblock[27][30] ),
    .S0(net50),
    .S1(net37),
    .X(_00807_));
 sky130_fd_sc_hd__mux4_2 _13990_ (.A0(\r1.regblock[28][30] ),
    .A1(\r1.regblock[29][30] ),
    .A2(\r1.regblock[30][30] ),
    .A3(\r1.regblock[31][30] ),
    .S0(net51),
    .S1(net37),
    .X(_00808_));
 sky130_fd_sc_hd__mux4_1 _13991_ (.A0(_00805_),
    .A1(_00806_),
    .A2(_00807_),
    .A3(_00808_),
    .S0(\c1.instruction1[22] ),
    .S1(\c1.instruction1[23] ),
    .X(_00809_));
 sky130_fd_sc_hd__mux4_1 _13992_ (.A0(\r1.regblock[0][29] ),
    .A1(\r1.regblock[1][29] ),
    .A2(\r1.regblock[2][29] ),
    .A3(\r1.regblock[3][29] ),
    .S0(net51),
    .S1(net37),
    .X(_00787_));
 sky130_fd_sc_hd__mux4_2 _13993_ (.A0(\r1.regblock[4][29] ),
    .A1(\r1.regblock[5][29] ),
    .A2(\r1.regblock[6][29] ),
    .A3(\r1.regblock[7][29] ),
    .S0(net51),
    .S1(net37),
    .X(_00788_));
 sky130_fd_sc_hd__mux4_1 _13994_ (.A0(\r1.regblock[8][29] ),
    .A1(\r1.regblock[9][29] ),
    .A2(\r1.regblock[10][29] ),
    .A3(\r1.regblock[11][29] ),
    .S0(net51),
    .S1(net37),
    .X(_00789_));
 sky130_fd_sc_hd__mux4_1 _13995_ (.A0(\r1.regblock[12][29] ),
    .A1(\r1.regblock[13][29] ),
    .A2(\r1.regblock[14][29] ),
    .A3(\r1.regblock[15][29] ),
    .S0(net51),
    .S1(net37),
    .X(_00790_));
 sky130_fd_sc_hd__mux4_2 _13996_ (.A0(_00787_),
    .A1(_00788_),
    .A2(_00789_),
    .A3(_00790_),
    .S0(net34),
    .S1(net32),
    .X(_00791_));
 sky130_fd_sc_hd__mux4_1 _13997_ (.A0(\r1.regblock[16][29] ),
    .A1(\r1.regblock[17][29] ),
    .A2(\r1.regblock[18][29] ),
    .A3(\r1.regblock[19][29] ),
    .S0(net51),
    .S1(net37),
    .X(_00792_));
 sky130_fd_sc_hd__mux4_2 _13998_ (.A0(\r1.regblock[20][29] ),
    .A1(\r1.regblock[21][29] ),
    .A2(\r1.regblock[22][29] ),
    .A3(\r1.regblock[23][29] ),
    .S0(net51),
    .S1(net37),
    .X(_00793_));
 sky130_fd_sc_hd__mux4_2 _13999_ (.A0(\r1.regblock[24][29] ),
    .A1(\r1.regblock[25][29] ),
    .A2(\r1.regblock[26][29] ),
    .A3(\r1.regblock[27][29] ),
    .S0(net50),
    .S1(net37),
    .X(_00794_));
 sky130_fd_sc_hd__mux4_2 _14000_ (.A0(\r1.regblock[28][29] ),
    .A1(\r1.regblock[29][29] ),
    .A2(\r1.regblock[30][29] ),
    .A3(\r1.regblock[31][29] ),
    .S0(net51),
    .S1(net37),
    .X(_00795_));
 sky130_fd_sc_hd__mux4_1 _14001_ (.A0(_00792_),
    .A1(_00793_),
    .A2(_00794_),
    .A3(_00795_),
    .S0(\c1.instruction1[22] ),
    .S1(\c1.instruction1[23] ),
    .X(_00796_));
 sky130_fd_sc_hd__mux4_1 _14002_ (.A0(\r1.regblock[0][28] ),
    .A1(\r1.regblock[1][28] ),
    .A2(\r1.regblock[2][28] ),
    .A3(\r1.regblock[3][28] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00774_));
 sky130_fd_sc_hd__mux4_2 _14003_ (.A0(\r1.regblock[4][28] ),
    .A1(\r1.regblock[5][28] ),
    .A2(\r1.regblock[6][28] ),
    .A3(\r1.regblock[7][28] ),
    .S0(net52),
    .S1(net36),
    .X(_00775_));
 sky130_fd_sc_hd__mux4_2 _14004_ (.A0(\r1.regblock[8][28] ),
    .A1(\r1.regblock[9][28] ),
    .A2(\r1.regblock[10][28] ),
    .A3(\r1.regblock[11][28] ),
    .S0(net52),
    .S1(net36),
    .X(_00776_));
 sky130_fd_sc_hd__mux4_1 _14005_ (.A0(\r1.regblock[12][28] ),
    .A1(\r1.regblock[13][28] ),
    .A2(\r1.regblock[14][28] ),
    .A3(\r1.regblock[15][28] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00777_));
 sky130_fd_sc_hd__mux4_2 _14006_ (.A0(_00774_),
    .A1(_00775_),
    .A2(_00776_),
    .A3(_00777_),
    .S0(net34),
    .S1(net32),
    .X(_00778_));
 sky130_fd_sc_hd__mux4_2 _14007_ (.A0(\r1.regblock[16][28] ),
    .A1(\r1.regblock[17][28] ),
    .A2(\r1.regblock[18][28] ),
    .A3(\r1.regblock[19][28] ),
    .S0(net51),
    .S1(net36),
    .X(_00779_));
 sky130_fd_sc_hd__mux4_1 _14008_ (.A0(\r1.regblock[20][28] ),
    .A1(\r1.regblock[21][28] ),
    .A2(\r1.regblock[22][28] ),
    .A3(\r1.regblock[23][28] ),
    .S0(net51),
    .S1(net36),
    .X(_00780_));
 sky130_fd_sc_hd__mux4_2 _14009_ (.A0(\r1.regblock[24][28] ),
    .A1(\r1.regblock[25][28] ),
    .A2(\r1.regblock[26][28] ),
    .A3(\r1.regblock[27][28] ),
    .S0(net51),
    .S1(net36),
    .X(_00781_));
 sky130_fd_sc_hd__mux4_2 _14010_ (.A0(\r1.regblock[28][28] ),
    .A1(\r1.regblock[29][28] ),
    .A2(\r1.regblock[30][28] ),
    .A3(\r1.regblock[31][28] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00782_));
 sky130_fd_sc_hd__mux4_1 _14011_ (.A0(_00779_),
    .A1(_00780_),
    .A2(_00781_),
    .A3(_00782_),
    .S0(net34),
    .S1(net32),
    .X(_00783_));
 sky130_fd_sc_hd__mux4_1 _14012_ (.A0(\r1.regblock[0][27] ),
    .A1(\r1.regblock[1][27] ),
    .A2(\r1.regblock[2][27] ),
    .A3(\r1.regblock[3][27] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00761_));
 sky130_fd_sc_hd__mux4_2 _14013_ (.A0(\r1.regblock[4][27] ),
    .A1(\r1.regblock[5][27] ),
    .A2(\r1.regblock[6][27] ),
    .A3(\r1.regblock[7][27] ),
    .S0(net52),
    .S1(net36),
    .X(_00762_));
 sky130_fd_sc_hd__mux4_2 _14014_ (.A0(\r1.regblock[8][27] ),
    .A1(\r1.regblock[9][27] ),
    .A2(\r1.regblock[10][27] ),
    .A3(\r1.regblock[11][27] ),
    .S0(net52),
    .S1(net36),
    .X(_00763_));
 sky130_fd_sc_hd__mux4_2 _14015_ (.A0(\r1.regblock[12][27] ),
    .A1(\r1.regblock[13][27] ),
    .A2(\r1.regblock[14][27] ),
    .A3(\r1.regblock[15][27] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00764_));
 sky130_fd_sc_hd__mux4_2 _14016_ (.A0(_00761_),
    .A1(_00762_),
    .A2(_00763_),
    .A3(_00764_),
    .S0(net34),
    .S1(net32),
    .X(_00765_));
 sky130_fd_sc_hd__mux4_2 _14017_ (.A0(\r1.regblock[16][27] ),
    .A1(\r1.regblock[17][27] ),
    .A2(\r1.regblock[18][27] ),
    .A3(\r1.regblock[19][27] ),
    .S0(net51),
    .S1(net36),
    .X(_00766_));
 sky130_fd_sc_hd__mux4_1 _14018_ (.A0(\r1.regblock[20][27] ),
    .A1(\r1.regblock[21][27] ),
    .A2(\r1.regblock[22][27] ),
    .A3(\r1.regblock[23][27] ),
    .S0(net51),
    .S1(net36),
    .X(_00767_));
 sky130_fd_sc_hd__mux4_1 _14019_ (.A0(\r1.regblock[24][27] ),
    .A1(\r1.regblock[25][27] ),
    .A2(\r1.regblock[26][27] ),
    .A3(\r1.regblock[27][27] ),
    .S0(net51),
    .S1(net36),
    .X(_00768_));
 sky130_fd_sc_hd__mux4_2 _14020_ (.A0(\r1.regblock[28][27] ),
    .A1(\r1.regblock[29][27] ),
    .A2(\r1.regblock[30][27] ),
    .A3(\r1.regblock[31][27] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00769_));
 sky130_fd_sc_hd__mux4_1 _14021_ (.A0(_00766_),
    .A1(_00767_),
    .A2(_00768_),
    .A3(_00769_),
    .S0(net34),
    .S1(net32),
    .X(_00770_));
 sky130_fd_sc_hd__mux4_1 _14022_ (.A0(\r1.regblock[0][26] ),
    .A1(\r1.regblock[1][26] ),
    .A2(\r1.regblock[2][26] ),
    .A3(\r1.regblock[3][26] ),
    .S0(net52),
    .S1(net36),
    .X(_00748_));
 sky130_fd_sc_hd__mux4_2 _14023_ (.A0(\r1.regblock[4][26] ),
    .A1(\r1.regblock[5][26] ),
    .A2(\r1.regblock[6][26] ),
    .A3(\r1.regblock[7][26] ),
    .S0(net52),
    .S1(net36),
    .X(_00749_));
 sky130_fd_sc_hd__mux4_2 _14024_ (.A0(\r1.regblock[8][26] ),
    .A1(\r1.regblock[9][26] ),
    .A2(\r1.regblock[10][26] ),
    .A3(\r1.regblock[11][26] ),
    .S0(net52),
    .S1(net36),
    .X(_00750_));
 sky130_fd_sc_hd__mux4_2 _14025_ (.A0(\r1.regblock[12][26] ),
    .A1(\r1.regblock[13][26] ),
    .A2(\r1.regblock[14][26] ),
    .A3(\r1.regblock[15][26] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00751_));
 sky130_fd_sc_hd__mux4_2 _14026_ (.A0(_00748_),
    .A1(_00749_),
    .A2(_00750_),
    .A3(_00751_),
    .S0(net34),
    .S1(net32),
    .X(_00752_));
 sky130_fd_sc_hd__mux4_2 _14027_ (.A0(\r1.regblock[16][26] ),
    .A1(\r1.regblock[17][26] ),
    .A2(\r1.regblock[18][26] ),
    .A3(\r1.regblock[19][26] ),
    .S0(net51),
    .S1(net36),
    .X(_00753_));
 sky130_fd_sc_hd__mux4_2 _14028_ (.A0(\r1.regblock[20][26] ),
    .A1(\r1.regblock[21][26] ),
    .A2(\r1.regblock[22][26] ),
    .A3(\r1.regblock[23][26] ),
    .S0(net51),
    .S1(net36),
    .X(_00754_));
 sky130_fd_sc_hd__mux4_1 _14029_ (.A0(\r1.regblock[24][26] ),
    .A1(\r1.regblock[25][26] ),
    .A2(\r1.regblock[26][26] ),
    .A3(\r1.regblock[27][26] ),
    .S0(net51),
    .S1(net36),
    .X(_00755_));
 sky130_fd_sc_hd__mux4_2 _14030_ (.A0(\r1.regblock[28][26] ),
    .A1(\r1.regblock[29][26] ),
    .A2(\r1.regblock[30][26] ),
    .A3(\r1.regblock[31][26] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00756_));
 sky130_fd_sc_hd__mux4_1 _14031_ (.A0(_00753_),
    .A1(_00754_),
    .A2(_00755_),
    .A3(_00756_),
    .S0(net34),
    .S1(net32),
    .X(_00757_));
 sky130_fd_sc_hd__mux4_1 _14032_ (.A0(\r1.regblock[0][25] ),
    .A1(\r1.regblock[1][25] ),
    .A2(\r1.regblock[2][25] ),
    .A3(\r1.regblock[3][25] ),
    .S0(net52),
    .S1(net36),
    .X(_00735_));
 sky130_fd_sc_hd__mux4_1 _14033_ (.A0(\r1.regblock[4][25] ),
    .A1(\r1.regblock[5][25] ),
    .A2(\r1.regblock[6][25] ),
    .A3(\r1.regblock[7][25] ),
    .S0(net52),
    .S1(net36),
    .X(_00736_));
 sky130_fd_sc_hd__mux4_2 _14034_ (.A0(\r1.regblock[8][25] ),
    .A1(\r1.regblock[9][25] ),
    .A2(\r1.regblock[10][25] ),
    .A3(\r1.regblock[11][25] ),
    .S0(net52),
    .S1(net38),
    .X(_00737_));
 sky130_fd_sc_hd__mux4_2 _14035_ (.A0(\r1.regblock[12][25] ),
    .A1(\r1.regblock[13][25] ),
    .A2(\r1.regblock[14][25] ),
    .A3(\r1.regblock[15][25] ),
    .S0(net52),
    .S1(net36),
    .X(_00738_));
 sky130_fd_sc_hd__mux4_2 _14036_ (.A0(_00735_),
    .A1(_00736_),
    .A2(_00737_),
    .A3(_00738_),
    .S0(net34),
    .S1(net32),
    .X(_00739_));
 sky130_fd_sc_hd__mux4_2 _14037_ (.A0(\r1.regblock[16][25] ),
    .A1(\r1.regblock[17][25] ),
    .A2(\r1.regblock[18][25] ),
    .A3(\r1.regblock[19][25] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00740_));
 sky130_fd_sc_hd__mux4_1 _14038_ (.A0(\r1.regblock[20][25] ),
    .A1(\r1.regblock[21][25] ),
    .A2(\r1.regblock[22][25] ),
    .A3(\r1.regblock[23][25] ),
    .S0(\c1.instruction1[20] ),
    .S1(net37),
    .X(_00741_));
 sky130_fd_sc_hd__mux4_2 _14039_ (.A0(\r1.regblock[24][25] ),
    .A1(\r1.regblock[25][25] ),
    .A2(\r1.regblock[26][25] ),
    .A3(\r1.regblock[27][25] ),
    .S0(\c1.instruction1[20] ),
    .S1(net37),
    .X(_00742_));
 sky130_fd_sc_hd__mux4_2 _14040_ (.A0(\r1.regblock[28][25] ),
    .A1(\r1.regblock[29][25] ),
    .A2(\r1.regblock[30][25] ),
    .A3(\r1.regblock[31][25] ),
    .S0(net51),
    .S1(net37),
    .X(_00743_));
 sky130_fd_sc_hd__mux4_1 _14041_ (.A0(_00740_),
    .A1(_00741_),
    .A2(_00742_),
    .A3(_00743_),
    .S0(net34),
    .S1(net32),
    .X(_00744_));
 sky130_fd_sc_hd__mux4_1 _14042_ (.A0(\r1.regblock[0][24] ),
    .A1(\r1.regblock[1][24] ),
    .A2(\r1.regblock[2][24] ),
    .A3(\r1.regblock[3][24] ),
    .S0(net52),
    .S1(net36),
    .X(_00722_));
 sky130_fd_sc_hd__mux4_2 _14043_ (.A0(\r1.regblock[4][24] ),
    .A1(\r1.regblock[5][24] ),
    .A2(\r1.regblock[6][24] ),
    .A3(\r1.regblock[7][24] ),
    .S0(net52),
    .S1(net36),
    .X(_00723_));
 sky130_fd_sc_hd__mux4_2 _14044_ (.A0(\r1.regblock[8][24] ),
    .A1(\r1.regblock[9][24] ),
    .A2(\r1.regblock[10][24] ),
    .A3(\r1.regblock[11][24] ),
    .S0(net43),
    .S1(net38),
    .X(_00724_));
 sky130_fd_sc_hd__mux4_1 _14045_ (.A0(\r1.regblock[12][24] ),
    .A1(\r1.regblock[13][24] ),
    .A2(\r1.regblock[14][24] ),
    .A3(\r1.regblock[15][24] ),
    .S0(net52),
    .S1(net36),
    .X(_00725_));
 sky130_fd_sc_hd__mux4_2 _14046_ (.A0(_00722_),
    .A1(_00723_),
    .A2(_00724_),
    .A3(_00725_),
    .S0(net34),
    .S1(net32),
    .X(_00726_));
 sky130_fd_sc_hd__mux4_2 _14047_ (.A0(\r1.regblock[16][24] ),
    .A1(\r1.regblock[17][24] ),
    .A2(\r1.regblock[18][24] ),
    .A3(\r1.regblock[19][24] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00727_));
 sky130_fd_sc_hd__mux4_2 _14048_ (.A0(\r1.regblock[20][24] ),
    .A1(\r1.regblock[21][24] ),
    .A2(\r1.regblock[22][24] ),
    .A3(\r1.regblock[23][24] ),
    .S0(\c1.instruction1[20] ),
    .S1(net37),
    .X(_00728_));
 sky130_fd_sc_hd__mux4_1 _14049_ (.A0(\r1.regblock[24][24] ),
    .A1(\r1.regblock[25][24] ),
    .A2(\r1.regblock[26][24] ),
    .A3(\r1.regblock[27][24] ),
    .S0(\c1.instruction1[20] ),
    .S1(net37),
    .X(_00729_));
 sky130_fd_sc_hd__mux4_1 _14050_ (.A0(\r1.regblock[28][24] ),
    .A1(\r1.regblock[29][24] ),
    .A2(\r1.regblock[30][24] ),
    .A3(\r1.regblock[31][24] ),
    .S0(\c1.instruction1[20] ),
    .S1(net37),
    .X(_00730_));
 sky130_fd_sc_hd__mux4_1 _14051_ (.A0(_00727_),
    .A1(_00728_),
    .A2(_00729_),
    .A3(_00730_),
    .S0(net34),
    .S1(net32),
    .X(_00731_));
 sky130_fd_sc_hd__mux4_1 _14052_ (.A0(\r1.regblock[0][23] ),
    .A1(\r1.regblock[1][23] ),
    .A2(\r1.regblock[2][23] ),
    .A3(\r1.regblock[3][23] ),
    .S0(net52),
    .S1(net36),
    .X(_00709_));
 sky130_fd_sc_hd__mux4_2 _14053_ (.A0(\r1.regblock[4][23] ),
    .A1(\r1.regblock[5][23] ),
    .A2(\r1.regblock[6][23] ),
    .A3(\r1.regblock[7][23] ),
    .S0(net52),
    .S1(net36),
    .X(_00710_));
 sky130_fd_sc_hd__mux4_2 _14054_ (.A0(\r1.regblock[8][23] ),
    .A1(\r1.regblock[9][23] ),
    .A2(\r1.regblock[10][23] ),
    .A3(\r1.regblock[11][23] ),
    .S0(net43),
    .S1(net38),
    .X(_00711_));
 sky130_fd_sc_hd__mux4_1 _14055_ (.A0(\r1.regblock[12][23] ),
    .A1(\r1.regblock[13][23] ),
    .A2(\r1.regblock[14][23] ),
    .A3(\r1.regblock[15][23] ),
    .S0(net52),
    .S1(net36),
    .X(_00712_));
 sky130_fd_sc_hd__mux4_2 _14056_ (.A0(_00709_),
    .A1(_00710_),
    .A2(_00711_),
    .A3(_00712_),
    .S0(net34),
    .S1(net32),
    .X(_00713_));
 sky130_fd_sc_hd__mux4_2 _14057_ (.A0(\r1.regblock[16][23] ),
    .A1(\r1.regblock[17][23] ),
    .A2(\r1.regblock[18][23] ),
    .A3(\r1.regblock[19][23] ),
    .S0(\c1.instruction1[20] ),
    .S1(net36),
    .X(_00714_));
 sky130_fd_sc_hd__mux4_2 _14058_ (.A0(\r1.regblock[20][23] ),
    .A1(\r1.regblock[21][23] ),
    .A2(\r1.regblock[22][23] ),
    .A3(\r1.regblock[23][23] ),
    .S0(\c1.instruction1[20] ),
    .S1(net37),
    .X(_00715_));
 sky130_fd_sc_hd__mux4_1 _14059_ (.A0(\r1.regblock[24][23] ),
    .A1(\r1.regblock[25][23] ),
    .A2(\r1.regblock[26][23] ),
    .A3(\r1.regblock[27][23] ),
    .S0(\c1.instruction1[20] ),
    .S1(net37),
    .X(_00716_));
 sky130_fd_sc_hd__mux4_2 _14060_ (.A0(\r1.regblock[28][23] ),
    .A1(\r1.regblock[29][23] ),
    .A2(\r1.regblock[30][23] ),
    .A3(\r1.regblock[31][23] ),
    .S0(net51),
    .S1(net37),
    .X(_00717_));
 sky130_fd_sc_hd__mux4_1 _14061_ (.A0(_00714_),
    .A1(_00715_),
    .A2(_00716_),
    .A3(_00717_),
    .S0(net34),
    .S1(net32),
    .X(_00718_));
 sky130_fd_sc_hd__mux4_1 _14062_ (.A0(\r1.regblock[0][22] ),
    .A1(\r1.regblock[1][22] ),
    .A2(\r1.regblock[2][22] ),
    .A3(\r1.regblock[3][22] ),
    .S0(net43),
    .S1(net38),
    .X(_00696_));
 sky130_fd_sc_hd__mux4_2 _14063_ (.A0(\r1.regblock[4][22] ),
    .A1(\r1.regblock[5][22] ),
    .A2(\r1.regblock[6][22] ),
    .A3(\r1.regblock[7][22] ),
    .S0(net43),
    .S1(net38),
    .X(_00697_));
 sky130_fd_sc_hd__mux4_2 _14064_ (.A0(\r1.regblock[8][22] ),
    .A1(\r1.regblock[9][22] ),
    .A2(\r1.regblock[10][22] ),
    .A3(\r1.regblock[11][22] ),
    .S0(net43),
    .S1(net38),
    .X(_00698_));
 sky130_fd_sc_hd__mux4_1 _14065_ (.A0(\r1.regblock[12][22] ),
    .A1(\r1.regblock[13][22] ),
    .A2(\r1.regblock[14][22] ),
    .A3(\r1.regblock[15][22] ),
    .S0(net43),
    .S1(net38),
    .X(_00699_));
 sky130_fd_sc_hd__mux4_2 _14066_ (.A0(_00696_),
    .A1(_00697_),
    .A2(_00698_),
    .A3(_00699_),
    .S0(net34),
    .S1(net32),
    .X(_00700_));
 sky130_fd_sc_hd__mux4_2 _14067_ (.A0(\r1.regblock[16][22] ),
    .A1(\r1.regblock[17][22] ),
    .A2(\r1.regblock[18][22] ),
    .A3(\r1.regblock[19][22] ),
    .S0(net43),
    .S1(net38),
    .X(_00701_));
 sky130_fd_sc_hd__mux4_2 _14068_ (.A0(\r1.regblock[20][22] ),
    .A1(\r1.regblock[21][22] ),
    .A2(\r1.regblock[22][22] ),
    .A3(\r1.regblock[23][22] ),
    .S0(net43),
    .S1(net38),
    .X(_00702_));
 sky130_fd_sc_hd__mux4_2 _14069_ (.A0(\r1.regblock[24][22] ),
    .A1(\r1.regblock[25][22] ),
    .A2(\r1.regblock[26][22] ),
    .A3(\r1.regblock[27][22] ),
    .S0(net43),
    .S1(net38),
    .X(_00703_));
 sky130_fd_sc_hd__mux4_1 _14070_ (.A0(\r1.regblock[28][22] ),
    .A1(\r1.regblock[29][22] ),
    .A2(\r1.regblock[30][22] ),
    .A3(\r1.regblock[31][22] ),
    .S0(net43),
    .S1(net38),
    .X(_00704_));
 sky130_fd_sc_hd__mux4_1 _14071_ (.A0(_00701_),
    .A1(_00702_),
    .A2(_00703_),
    .A3(_00704_),
    .S0(net34),
    .S1(net32),
    .X(_00705_));
 sky130_fd_sc_hd__mux4_1 _14072_ (.A0(\r1.regblock[0][21] ),
    .A1(\r1.regblock[1][21] ),
    .A2(\r1.regblock[2][21] ),
    .A3(\r1.regblock[3][21] ),
    .S0(net43),
    .S1(net38),
    .X(_00683_));
 sky130_fd_sc_hd__mux4_2 _14073_ (.A0(\r1.regblock[4][21] ),
    .A1(\r1.regblock[5][21] ),
    .A2(\r1.regblock[6][21] ),
    .A3(\r1.regblock[7][21] ),
    .S0(net43),
    .S1(net38),
    .X(_00684_));
 sky130_fd_sc_hd__mux4_2 _14074_ (.A0(\r1.regblock[8][21] ),
    .A1(\r1.regblock[9][21] ),
    .A2(\r1.regblock[10][21] ),
    .A3(\r1.regblock[11][21] ),
    .S0(net43),
    .S1(net38),
    .X(_00685_));
 sky130_fd_sc_hd__mux4_1 _14075_ (.A0(\r1.regblock[12][21] ),
    .A1(\r1.regblock[13][21] ),
    .A2(\r1.regblock[14][21] ),
    .A3(\r1.regblock[15][21] ),
    .S0(net43),
    .S1(net38),
    .X(_00686_));
 sky130_fd_sc_hd__mux4_2 _14076_ (.A0(_00683_),
    .A1(_00684_),
    .A2(_00685_),
    .A3(_00686_),
    .S0(net34),
    .S1(net32),
    .X(_00687_));
 sky130_fd_sc_hd__mux4_2 _14077_ (.A0(\r1.regblock[16][21] ),
    .A1(\r1.regblock[17][21] ),
    .A2(\r1.regblock[18][21] ),
    .A3(\r1.regblock[19][21] ),
    .S0(net43),
    .S1(net38),
    .X(_00688_));
 sky130_fd_sc_hd__mux4_1 _14078_ (.A0(\r1.regblock[20][21] ),
    .A1(\r1.regblock[21][21] ),
    .A2(\r1.regblock[22][21] ),
    .A3(\r1.regblock[23][21] ),
    .S0(net43),
    .S1(net38),
    .X(_00689_));
 sky130_fd_sc_hd__mux4_2 _14079_ (.A0(\r1.regblock[24][21] ),
    .A1(\r1.regblock[25][21] ),
    .A2(\r1.regblock[26][21] ),
    .A3(\r1.regblock[27][21] ),
    .S0(net43),
    .S1(net38),
    .X(_00690_));
 sky130_fd_sc_hd__mux4_1 _14080_ (.A0(\r1.regblock[28][21] ),
    .A1(\r1.regblock[29][21] ),
    .A2(\r1.regblock[30][21] ),
    .A3(\r1.regblock[31][21] ),
    .S0(net43),
    .S1(net38),
    .X(_00691_));
 sky130_fd_sc_hd__mux4_1 _14081_ (.A0(_00688_),
    .A1(_00689_),
    .A2(_00690_),
    .A3(_00691_),
    .S0(net34),
    .S1(net32),
    .X(_00692_));
 sky130_fd_sc_hd__mux4_1 _14082_ (.A0(\r1.regblock[0][20] ),
    .A1(\r1.regblock[1][20] ),
    .A2(\r1.regblock[2][20] ),
    .A3(\r1.regblock[3][20] ),
    .S0(net43),
    .S1(net38),
    .X(_00670_));
 sky130_fd_sc_hd__mux4_2 _14083_ (.A0(\r1.regblock[4][20] ),
    .A1(\r1.regblock[5][20] ),
    .A2(\r1.regblock[6][20] ),
    .A3(\r1.regblock[7][20] ),
    .S0(net43),
    .S1(net38),
    .X(_00671_));
 sky130_fd_sc_hd__mux4_1 _14084_ (.A0(\r1.regblock[8][20] ),
    .A1(\r1.regblock[9][20] ),
    .A2(\r1.regblock[10][20] ),
    .A3(\r1.regblock[11][20] ),
    .S0(net43),
    .S1(net38),
    .X(_00672_));
 sky130_fd_sc_hd__mux4_1 _14085_ (.A0(\r1.regblock[12][20] ),
    .A1(\r1.regblock[13][20] ),
    .A2(\r1.regblock[14][20] ),
    .A3(\r1.regblock[15][20] ),
    .S0(net43),
    .S1(net38),
    .X(_00673_));
 sky130_fd_sc_hd__mux4_2 _14086_ (.A0(_00670_),
    .A1(_00671_),
    .A2(_00672_),
    .A3(_00673_),
    .S0(net34),
    .S1(net32),
    .X(_00674_));
 sky130_fd_sc_hd__mux4_2 _14087_ (.A0(\r1.regblock[16][20] ),
    .A1(\r1.regblock[17][20] ),
    .A2(\r1.regblock[18][20] ),
    .A3(\r1.regblock[19][20] ),
    .S0(net43),
    .S1(net38),
    .X(_00675_));
 sky130_fd_sc_hd__mux4_2 _14088_ (.A0(\r1.regblock[20][20] ),
    .A1(\r1.regblock[21][20] ),
    .A2(\r1.regblock[22][20] ),
    .A3(\r1.regblock[23][20] ),
    .S0(net43),
    .S1(net38),
    .X(_00676_));
 sky130_fd_sc_hd__mux4_1 _14089_ (.A0(\r1.regblock[24][20] ),
    .A1(\r1.regblock[25][20] ),
    .A2(\r1.regblock[26][20] ),
    .A3(\r1.regblock[27][20] ),
    .S0(net43),
    .S1(net38),
    .X(_00677_));
 sky130_fd_sc_hd__mux4_1 _14090_ (.A0(\r1.regblock[28][20] ),
    .A1(\r1.regblock[29][20] ),
    .A2(\r1.regblock[30][20] ),
    .A3(\r1.regblock[31][20] ),
    .S0(net43),
    .S1(net38),
    .X(_00678_));
 sky130_fd_sc_hd__mux4_1 _14091_ (.A0(_00675_),
    .A1(_00676_),
    .A2(_00677_),
    .A3(_00678_),
    .S0(net34),
    .S1(net32),
    .X(_00679_));
 sky130_fd_sc_hd__mux4_1 _14092_ (.A0(\r1.regblock[0][19] ),
    .A1(\r1.regblock[1][19] ),
    .A2(\r1.regblock[2][19] ),
    .A3(\r1.regblock[3][19] ),
    .S0(net45),
    .S1(net41),
    .X(_00657_));
 sky130_fd_sc_hd__mux4_2 _14093_ (.A0(\r1.regblock[4][19] ),
    .A1(\r1.regblock[5][19] ),
    .A2(\r1.regblock[6][19] ),
    .A3(\r1.regblock[7][19] ),
    .S0(net46),
    .S1(net42),
    .X(_00658_));
 sky130_fd_sc_hd__mux4_1 _14094_ (.A0(\r1.regblock[8][19] ),
    .A1(\r1.regblock[9][19] ),
    .A2(\r1.regblock[10][19] ),
    .A3(\r1.regblock[11][19] ),
    .S0(net46),
    .S1(net41),
    .X(_00659_));
 sky130_fd_sc_hd__mux4_1 _14095_ (.A0(\r1.regblock[12][19] ),
    .A1(\r1.regblock[13][19] ),
    .A2(\r1.regblock[14][19] ),
    .A3(\r1.regblock[15][19] ),
    .S0(net45),
    .S1(net41),
    .X(_00660_));
 sky130_fd_sc_hd__mux4_2 _14096_ (.A0(_00657_),
    .A1(_00658_),
    .A2(_00659_),
    .A3(_00660_),
    .S0(net35),
    .S1(net33),
    .X(_00661_));
 sky130_fd_sc_hd__mux4_2 _14097_ (.A0(\r1.regblock[16][19] ),
    .A1(\r1.regblock[17][19] ),
    .A2(\r1.regblock[18][19] ),
    .A3(\r1.regblock[19][19] ),
    .S0(net45),
    .S1(net41),
    .X(_00662_));
 sky130_fd_sc_hd__mux4_1 _14098_ (.A0(\r1.regblock[20][19] ),
    .A1(\r1.regblock[21][19] ),
    .A2(\r1.regblock[22][19] ),
    .A3(\r1.regblock[23][19] ),
    .S0(net45),
    .S1(net41),
    .X(_00663_));
 sky130_fd_sc_hd__mux4_2 _14099_ (.A0(\r1.regblock[24][19] ),
    .A1(\r1.regblock[25][19] ),
    .A2(\r1.regblock[26][19] ),
    .A3(\r1.regblock[27][19] ),
    .S0(net45),
    .S1(net41),
    .X(_00664_));
 sky130_fd_sc_hd__mux4_2 _14100_ (.A0(\r1.regblock[28][19] ),
    .A1(\r1.regblock[29][19] ),
    .A2(\r1.regblock[30][19] ),
    .A3(\r1.regblock[31][19] ),
    .S0(net45),
    .S1(net41),
    .X(_00665_));
 sky130_fd_sc_hd__mux4_1 _14101_ (.A0(_00662_),
    .A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00666_));
 sky130_fd_sc_hd__mux4_1 _14102_ (.A0(\r1.regblock[0][18] ),
    .A1(\r1.regblock[1][18] ),
    .A2(\r1.regblock[2][18] ),
    .A3(\r1.regblock[3][18] ),
    .S0(net45),
    .S1(net41),
    .X(_00644_));
 sky130_fd_sc_hd__mux4_2 _14103_ (.A0(\r1.regblock[4][18] ),
    .A1(\r1.regblock[5][18] ),
    .A2(\r1.regblock[6][18] ),
    .A3(\r1.regblock[7][18] ),
    .S0(net46),
    .S1(net42),
    .X(_00645_));
 sky130_fd_sc_hd__mux4_1 _14104_ (.A0(\r1.regblock[8][18] ),
    .A1(\r1.regblock[9][18] ),
    .A2(\r1.regblock[10][18] ),
    .A3(\r1.regblock[11][18] ),
    .S0(net45),
    .S1(net41),
    .X(_00646_));
 sky130_fd_sc_hd__mux4_1 _14105_ (.A0(\r1.regblock[12][18] ),
    .A1(\r1.regblock[13][18] ),
    .A2(\r1.regblock[14][18] ),
    .A3(\r1.regblock[15][18] ),
    .S0(net45),
    .S1(net41),
    .X(_00647_));
 sky130_fd_sc_hd__mux4_2 _14106_ (.A0(_00644_),
    .A1(_00645_),
    .A2(_00646_),
    .A3(_00647_),
    .S0(net35),
    .S1(net33),
    .X(_00648_));
 sky130_fd_sc_hd__mux4_2 _14107_ (.A0(\r1.regblock[16][18] ),
    .A1(\r1.regblock[17][18] ),
    .A2(\r1.regblock[18][18] ),
    .A3(\r1.regblock[19][18] ),
    .S0(net45),
    .S1(net41),
    .X(_00649_));
 sky130_fd_sc_hd__mux4_1 _14108_ (.A0(\r1.regblock[20][18] ),
    .A1(\r1.regblock[21][18] ),
    .A2(\r1.regblock[22][18] ),
    .A3(\r1.regblock[23][18] ),
    .S0(net45),
    .S1(net41),
    .X(_00650_));
 sky130_fd_sc_hd__mux4_2 _14109_ (.A0(\r1.regblock[24][18] ),
    .A1(\r1.regblock[25][18] ),
    .A2(\r1.regblock[26][18] ),
    .A3(\r1.regblock[27][18] ),
    .S0(net45),
    .S1(net41),
    .X(_00651_));
 sky130_fd_sc_hd__mux4_2 _14110_ (.A0(\r1.regblock[28][18] ),
    .A1(\r1.regblock[29][18] ),
    .A2(\r1.regblock[30][18] ),
    .A3(\r1.regblock[31][18] ),
    .S0(net45),
    .S1(net41),
    .X(_00652_));
 sky130_fd_sc_hd__mux4_1 _14111_ (.A0(_00649_),
    .A1(_00650_),
    .A2(_00651_),
    .A3(_00652_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00653_));
 sky130_fd_sc_hd__mux4_1 _14112_ (.A0(\r1.regblock[0][17] ),
    .A1(\r1.regblock[1][17] ),
    .A2(\r1.regblock[2][17] ),
    .A3(\r1.regblock[3][17] ),
    .S0(net45),
    .S1(net41),
    .X(_00631_));
 sky130_fd_sc_hd__mux4_2 _14113_ (.A0(\r1.regblock[4][17] ),
    .A1(\r1.regblock[5][17] ),
    .A2(\r1.regblock[6][17] ),
    .A3(\r1.regblock[7][17] ),
    .S0(net46),
    .S1(net42),
    .X(_00632_));
 sky130_fd_sc_hd__mux4_1 _14114_ (.A0(\r1.regblock[8][17] ),
    .A1(\r1.regblock[9][17] ),
    .A2(\r1.regblock[10][17] ),
    .A3(\r1.regblock[11][17] ),
    .S0(net45),
    .S1(net41),
    .X(_00633_));
 sky130_fd_sc_hd__mux4_1 _14115_ (.A0(\r1.regblock[12][17] ),
    .A1(\r1.regblock[13][17] ),
    .A2(\r1.regblock[14][17] ),
    .A3(\r1.regblock[15][17] ),
    .S0(net45),
    .S1(net41),
    .X(_00634_));
 sky130_fd_sc_hd__mux4_2 _14116_ (.A0(_00631_),
    .A1(_00632_),
    .A2(_00633_),
    .A3(_00634_),
    .S0(net35),
    .S1(net33),
    .X(_00635_));
 sky130_fd_sc_hd__mux4_2 _14117_ (.A0(\r1.regblock[16][17] ),
    .A1(\r1.regblock[17][17] ),
    .A2(\r1.regblock[18][17] ),
    .A3(\r1.regblock[19][17] ),
    .S0(net45),
    .S1(net41),
    .X(_00636_));
 sky130_fd_sc_hd__mux4_1 _14118_ (.A0(\r1.regblock[20][17] ),
    .A1(\r1.regblock[21][17] ),
    .A2(\r1.regblock[22][17] ),
    .A3(\r1.regblock[23][17] ),
    .S0(net45),
    .S1(net41),
    .X(_00637_));
 sky130_fd_sc_hd__mux4_2 _14119_ (.A0(\r1.regblock[24][17] ),
    .A1(\r1.regblock[25][17] ),
    .A2(\r1.regblock[26][17] ),
    .A3(\r1.regblock[27][17] ),
    .S0(net45),
    .S1(net41),
    .X(_00638_));
 sky130_fd_sc_hd__mux4_2 _14120_ (.A0(\r1.regblock[28][17] ),
    .A1(\r1.regblock[29][17] ),
    .A2(\r1.regblock[30][17] ),
    .A3(\r1.regblock[31][17] ),
    .S0(net45),
    .S1(net41),
    .X(_00639_));
 sky130_fd_sc_hd__mux4_1 _14121_ (.A0(_00636_),
    .A1(_00637_),
    .A2(_00638_),
    .A3(_00639_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00640_));
 sky130_fd_sc_hd__mux4_2 _14122_ (.A0(\r1.regblock[0][16] ),
    .A1(\r1.regblock[1][16] ),
    .A2(\r1.regblock[2][16] ),
    .A3(\r1.regblock[3][16] ),
    .S0(net45),
    .S1(net41),
    .X(_00618_));
 sky130_fd_sc_hd__mux4_2 _14123_ (.A0(\r1.regblock[4][16] ),
    .A1(\r1.regblock[5][16] ),
    .A2(\r1.regblock[6][16] ),
    .A3(\r1.regblock[7][16] ),
    .S0(net46),
    .S1(net42),
    .X(_00619_));
 sky130_fd_sc_hd__mux4_1 _14124_ (.A0(\r1.regblock[8][16] ),
    .A1(\r1.regblock[9][16] ),
    .A2(\r1.regblock[10][16] ),
    .A3(\r1.regblock[11][16] ),
    .S0(net45),
    .S1(net41),
    .X(_00620_));
 sky130_fd_sc_hd__mux4_1 _14125_ (.A0(\r1.regblock[12][16] ),
    .A1(\r1.regblock[13][16] ),
    .A2(\r1.regblock[14][16] ),
    .A3(\r1.regblock[15][16] ),
    .S0(net45),
    .S1(net41),
    .X(_00621_));
 sky130_fd_sc_hd__mux4_2 _14126_ (.A0(_00618_),
    .A1(_00619_),
    .A2(_00620_),
    .A3(_00621_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00622_));
 sky130_fd_sc_hd__mux4_2 _14127_ (.A0(\r1.regblock[16][16] ),
    .A1(\r1.regblock[17][16] ),
    .A2(\r1.regblock[18][16] ),
    .A3(\r1.regblock[19][16] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00623_));
 sky130_fd_sc_hd__mux4_2 _14128_ (.A0(\r1.regblock[20][16] ),
    .A1(\r1.regblock[21][16] ),
    .A2(\r1.regblock[22][16] ),
    .A3(\r1.regblock[23][16] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00624_));
 sky130_fd_sc_hd__mux4_2 _14129_ (.A0(\r1.regblock[24][16] ),
    .A1(\r1.regblock[25][16] ),
    .A2(\r1.regblock[26][16] ),
    .A3(\r1.regblock[27][16] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00625_));
 sky130_fd_sc_hd__mux4_1 _14130_ (.A0(\r1.regblock[28][16] ),
    .A1(\r1.regblock[29][16] ),
    .A2(\r1.regblock[30][16] ),
    .A3(\r1.regblock[31][16] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00626_));
 sky130_fd_sc_hd__mux4_2 _14131_ (.A0(_00623_),
    .A1(_00624_),
    .A2(_00625_),
    .A3(_00626_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00627_));
 sky130_fd_sc_hd__mux4_1 _14132_ (.A0(\r1.regblock[0][15] ),
    .A1(\r1.regblock[1][15] ),
    .A2(\r1.regblock[2][15] ),
    .A3(\r1.regblock[3][15] ),
    .S0(net45),
    .S1(net41),
    .X(_00605_));
 sky130_fd_sc_hd__mux4_2 _14133_ (.A0(\r1.regblock[4][15] ),
    .A1(\r1.regblock[5][15] ),
    .A2(\r1.regblock[6][15] ),
    .A3(\r1.regblock[7][15] ),
    .S0(net46),
    .S1(net42),
    .X(_00606_));
 sky130_fd_sc_hd__mux4_1 _14134_ (.A0(\r1.regblock[8][15] ),
    .A1(\r1.regblock[9][15] ),
    .A2(\r1.regblock[10][15] ),
    .A3(\r1.regblock[11][15] ),
    .S0(net45),
    .S1(net41),
    .X(_00607_));
 sky130_fd_sc_hd__mux4_2 _14135_ (.A0(\r1.regblock[12][15] ),
    .A1(\r1.regblock[13][15] ),
    .A2(\r1.regblock[14][15] ),
    .A3(\r1.regblock[15][15] ),
    .S0(net45),
    .S1(net41),
    .X(_00608_));
 sky130_fd_sc_hd__mux4_2 _14136_ (.A0(_00605_),
    .A1(_00606_),
    .A2(_00607_),
    .A3(_00608_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00609_));
 sky130_fd_sc_hd__mux4_1 _14137_ (.A0(\r1.regblock[16][15] ),
    .A1(\r1.regblock[17][15] ),
    .A2(\r1.regblock[18][15] ),
    .A3(\r1.regblock[19][15] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00610_));
 sky130_fd_sc_hd__mux4_2 _14138_ (.A0(\r1.regblock[20][15] ),
    .A1(\r1.regblock[21][15] ),
    .A2(\r1.regblock[22][15] ),
    .A3(\r1.regblock[23][15] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00611_));
 sky130_fd_sc_hd__mux4_2 _14139_ (.A0(\r1.regblock[24][15] ),
    .A1(\r1.regblock[25][15] ),
    .A2(\r1.regblock[26][15] ),
    .A3(\r1.regblock[27][15] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00612_));
 sky130_fd_sc_hd__mux4_1 _14140_ (.A0(\r1.regblock[28][15] ),
    .A1(\r1.regblock[29][15] ),
    .A2(\r1.regblock[30][15] ),
    .A3(\r1.regblock[31][15] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00613_));
 sky130_fd_sc_hd__mux4_1 _14141_ (.A0(_00610_),
    .A1(_00611_),
    .A2(_00612_),
    .A3(_00613_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00614_));
 sky130_fd_sc_hd__mux4_1 _14142_ (.A0(\r1.regblock[0][14] ),
    .A1(\r1.regblock[1][14] ),
    .A2(\r1.regblock[2][14] ),
    .A3(\r1.regblock[3][14] ),
    .S0(net45),
    .S1(net41),
    .X(_00592_));
 sky130_fd_sc_hd__mux4_2 _14143_ (.A0(\r1.regblock[4][14] ),
    .A1(\r1.regblock[5][14] ),
    .A2(\r1.regblock[6][14] ),
    .A3(\r1.regblock[7][14] ),
    .S0(net46),
    .S1(net42),
    .X(_00593_));
 sky130_fd_sc_hd__mux4_1 _14144_ (.A0(\r1.regblock[8][14] ),
    .A1(\r1.regblock[9][14] ),
    .A2(\r1.regblock[10][14] ),
    .A3(\r1.regblock[11][14] ),
    .S0(net45),
    .S1(net41),
    .X(_00594_));
 sky130_fd_sc_hd__mux4_2 _14145_ (.A0(\r1.regblock[12][14] ),
    .A1(\r1.regblock[13][14] ),
    .A2(\r1.regblock[14][14] ),
    .A3(\r1.regblock[15][14] ),
    .S0(net45),
    .S1(net41),
    .X(_00595_));
 sky130_fd_sc_hd__mux4_2 _14146_ (.A0(_00592_),
    .A1(_00593_),
    .A2(_00594_),
    .A3(_00595_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00596_));
 sky130_fd_sc_hd__mux4_1 _14147_ (.A0(\r1.regblock[16][14] ),
    .A1(\r1.regblock[17][14] ),
    .A2(\r1.regblock[18][14] ),
    .A3(\r1.regblock[19][14] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00597_));
 sky130_fd_sc_hd__mux4_2 _14148_ (.A0(\r1.regblock[20][14] ),
    .A1(\r1.regblock[21][14] ),
    .A2(\r1.regblock[22][14] ),
    .A3(\r1.regblock[23][14] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00598_));
 sky130_fd_sc_hd__mux4_1 _14149_ (.A0(\r1.regblock[24][14] ),
    .A1(\r1.regblock[25][14] ),
    .A2(\r1.regblock[26][14] ),
    .A3(\r1.regblock[27][14] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00599_));
 sky130_fd_sc_hd__mux4_1 _14150_ (.A0(\r1.regblock[28][14] ),
    .A1(\r1.regblock[29][14] ),
    .A2(\r1.regblock[30][14] ),
    .A3(\r1.regblock[31][14] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00600_));
 sky130_fd_sc_hd__mux4_1 _14151_ (.A0(_00597_),
    .A1(_00598_),
    .A2(_00599_),
    .A3(_00600_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00601_));
 sky130_fd_sc_hd__mux4_1 _14152_ (.A0(\r1.regblock[0][13] ),
    .A1(\r1.regblock[1][13] ),
    .A2(\r1.regblock[2][13] ),
    .A3(\r1.regblock[3][13] ),
    .S0(net44),
    .S1(net42),
    .X(_00579_));
 sky130_fd_sc_hd__mux4_2 _14153_ (.A0(\r1.regblock[4][13] ),
    .A1(\r1.regblock[5][13] ),
    .A2(\r1.regblock[6][13] ),
    .A3(\r1.regblock[7][13] ),
    .S0(net46),
    .S1(net42),
    .X(_00580_));
 sky130_fd_sc_hd__mux4_1 _14154_ (.A0(\r1.regblock[8][13] ),
    .A1(\r1.regblock[9][13] ),
    .A2(\r1.regblock[10][13] ),
    .A3(\r1.regblock[11][13] ),
    .S0(net44),
    .S1(net42),
    .X(_00581_));
 sky130_fd_sc_hd__mux4_2 _14155_ (.A0(\r1.regblock[12][13] ),
    .A1(\r1.regblock[13][13] ),
    .A2(\r1.regblock[14][13] ),
    .A3(\r1.regblock[15][13] ),
    .S0(net46),
    .S1(net42),
    .X(_00582_));
 sky130_fd_sc_hd__mux4_2 _14156_ (.A0(_00579_),
    .A1(_00580_),
    .A2(_00581_),
    .A3(_00582_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00583_));
 sky130_fd_sc_hd__mux4_2 _14157_ (.A0(\r1.regblock[16][13] ),
    .A1(\r1.regblock[17][13] ),
    .A2(\r1.regblock[18][13] ),
    .A3(\r1.regblock[19][13] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00584_));
 sky130_fd_sc_hd__mux4_2 _14158_ (.A0(\r1.regblock[20][13] ),
    .A1(\r1.regblock[21][13] ),
    .A2(\r1.regblock[22][13] ),
    .A3(\r1.regblock[23][13] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00585_));
 sky130_fd_sc_hd__mux4_1 _14159_ (.A0(\r1.regblock[24][13] ),
    .A1(\r1.regblock[25][13] ),
    .A2(\r1.regblock[26][13] ),
    .A3(\r1.regblock[27][13] ),
    .S0(net44),
    .S1(net42),
    .X(_00586_));
 sky130_fd_sc_hd__mux4_2 _14160_ (.A0(\r1.regblock[28][13] ),
    .A1(\r1.regblock[29][13] ),
    .A2(\r1.regblock[30][13] ),
    .A3(\r1.regblock[31][13] ),
    .S0(net44),
    .S1(net42),
    .X(_00587_));
 sky130_fd_sc_hd__mux4_1 _14161_ (.A0(_00584_),
    .A1(_00585_),
    .A2(_00586_),
    .A3(_00587_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00588_));
 sky130_fd_sc_hd__mux4_2 _14162_ (.A0(\r1.regblock[0][12] ),
    .A1(\r1.regblock[1][12] ),
    .A2(\r1.regblock[2][12] ),
    .A3(\r1.regblock[3][12] ),
    .S0(net44),
    .S1(net42),
    .X(_00566_));
 sky130_fd_sc_hd__mux4_2 _14163_ (.A0(\r1.regblock[4][12] ),
    .A1(\r1.regblock[5][12] ),
    .A2(\r1.regblock[6][12] ),
    .A3(\r1.regblock[7][12] ),
    .S0(net46),
    .S1(net42),
    .X(_00567_));
 sky130_fd_sc_hd__mux4_1 _14164_ (.A0(\r1.regblock[8][12] ),
    .A1(\r1.regblock[9][12] ),
    .A2(\r1.regblock[10][12] ),
    .A3(\r1.regblock[11][12] ),
    .S0(net44),
    .S1(net42),
    .X(_00568_));
 sky130_fd_sc_hd__mux4_2 _14165_ (.A0(\r1.regblock[12][12] ),
    .A1(\r1.regblock[13][12] ),
    .A2(\r1.regblock[14][12] ),
    .A3(\r1.regblock[15][12] ),
    .S0(net46),
    .S1(net42),
    .X(_00569_));
 sky130_fd_sc_hd__mux4_2 _14166_ (.A0(_00566_),
    .A1(_00567_),
    .A2(_00568_),
    .A3(_00569_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00570_));
 sky130_fd_sc_hd__mux4_2 _14167_ (.A0(\r1.regblock[16][12] ),
    .A1(\r1.regblock[17][12] ),
    .A2(\r1.regblock[18][12] ),
    .A3(\r1.regblock[19][12] ),
    .S0(net44),
    .S1(\c1.instruction1[21] ),
    .X(_00571_));
 sky130_fd_sc_hd__mux4_2 _14168_ (.A0(\r1.regblock[20][12] ),
    .A1(\r1.regblock[21][12] ),
    .A2(\r1.regblock[22][12] ),
    .A3(\r1.regblock[23][12] ),
    .S0(net44),
    .S1(net42),
    .X(_00572_));
 sky130_fd_sc_hd__mux4_1 _14169_ (.A0(\r1.regblock[24][12] ),
    .A1(\r1.regblock[25][12] ),
    .A2(\r1.regblock[26][12] ),
    .A3(\r1.regblock[27][12] ),
    .S0(net44),
    .S1(net42),
    .X(_00573_));
 sky130_fd_sc_hd__mux4_1 _14170_ (.A0(\r1.regblock[28][12] ),
    .A1(\r1.regblock[29][12] ),
    .A2(\r1.regblock[30][12] ),
    .A3(\r1.regblock[31][12] ),
    .S0(net44),
    .S1(net42),
    .X(_00574_));
 sky130_fd_sc_hd__mux4_1 _14171_ (.A0(_00571_),
    .A1(_00572_),
    .A2(_00573_),
    .A3(_00574_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00575_));
 sky130_fd_sc_hd__mux4_2 _14172_ (.A0(\r1.regblock[0][11] ),
    .A1(\r1.regblock[1][11] ),
    .A2(\r1.regblock[2][11] ),
    .A3(\r1.regblock[3][11] ),
    .S0(net44),
    .S1(net42),
    .X(_00553_));
 sky130_fd_sc_hd__mux4_2 _14173_ (.A0(\r1.regblock[4][11] ),
    .A1(\r1.regblock[5][11] ),
    .A2(\r1.regblock[6][11] ),
    .A3(\r1.regblock[7][11] ),
    .S0(net46),
    .S1(net42),
    .X(_00554_));
 sky130_fd_sc_hd__mux4_1 _14174_ (.A0(\r1.regblock[8][11] ),
    .A1(\r1.regblock[9][11] ),
    .A2(\r1.regblock[10][11] ),
    .A3(\r1.regblock[11][11] ),
    .S0(net46),
    .S1(net42),
    .X(_00555_));
 sky130_fd_sc_hd__mux4_1 _14175_ (.A0(\r1.regblock[12][11] ),
    .A1(\r1.regblock[13][11] ),
    .A2(\r1.regblock[14][11] ),
    .A3(\r1.regblock[15][11] ),
    .S0(net46),
    .S1(net42),
    .X(_00556_));
 sky130_fd_sc_hd__mux4_2 _14176_ (.A0(_00553_),
    .A1(_00554_),
    .A2(_00555_),
    .A3(_00556_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00557_));
 sky130_fd_sc_hd__mux4_2 _14177_ (.A0(\r1.regblock[16][11] ),
    .A1(\r1.regblock[17][11] ),
    .A2(\r1.regblock[18][11] ),
    .A3(\r1.regblock[19][11] ),
    .S0(net44),
    .S1(net42),
    .X(_00558_));
 sky130_fd_sc_hd__mux4_2 _14178_ (.A0(\r1.regblock[20][11] ),
    .A1(\r1.regblock[21][11] ),
    .A2(\r1.regblock[22][11] ),
    .A3(\r1.regblock[23][11] ),
    .S0(net44),
    .S1(net42),
    .X(_00559_));
 sky130_fd_sc_hd__mux4_2 _14179_ (.A0(\r1.regblock[24][11] ),
    .A1(\r1.regblock[25][11] ),
    .A2(\r1.regblock[26][11] ),
    .A3(\r1.regblock[27][11] ),
    .S0(net44),
    .S1(net42),
    .X(_00560_));
 sky130_fd_sc_hd__mux4_2 _14180_ (.A0(\r1.regblock[28][11] ),
    .A1(\r1.regblock[29][11] ),
    .A2(\r1.regblock[30][11] ),
    .A3(\r1.regblock[31][11] ),
    .S0(net44),
    .S1(net42),
    .X(_00561_));
 sky130_fd_sc_hd__mux4_1 _14181_ (.A0(_00558_),
    .A1(_00559_),
    .A2(_00560_),
    .A3(_00561_),
    .S0(\c1.instruction1[22] ),
    .S1(net33),
    .X(_00562_));
 sky130_fd_sc_hd__mux4_1 _14182_ (.A0(\r1.regblock[0][10] ),
    .A1(\r1.regblock[1][10] ),
    .A2(\r1.regblock[2][10] ),
    .A3(\r1.regblock[3][10] ),
    .S0(net48),
    .S1(net39),
    .X(_00540_));
 sky130_fd_sc_hd__mux4_2 _14183_ (.A0(\r1.regblock[4][10] ),
    .A1(\r1.regblock[5][10] ),
    .A2(\r1.regblock[6][10] ),
    .A3(\r1.regblock[7][10] ),
    .S0(net48),
    .S1(net39),
    .X(_00541_));
 sky130_fd_sc_hd__mux4_1 _14184_ (.A0(\r1.regblock[8][10] ),
    .A1(\r1.regblock[9][10] ),
    .A2(\r1.regblock[10][10] ),
    .A3(\r1.regblock[11][10] ),
    .S0(net48),
    .S1(net39),
    .X(_00542_));
 sky130_fd_sc_hd__mux4_1 _14185_ (.A0(\r1.regblock[12][10] ),
    .A1(\r1.regblock[13][10] ),
    .A2(\r1.regblock[14][10] ),
    .A3(\r1.regblock[15][10] ),
    .S0(net48),
    .S1(net39),
    .X(_00543_));
 sky130_fd_sc_hd__mux4_2 _14186_ (.A0(_00540_),
    .A1(_00541_),
    .A2(_00542_),
    .A3(_00543_),
    .S0(net35),
    .S1(net33),
    .X(_00544_));
 sky130_fd_sc_hd__mux4_2 _14187_ (.A0(\r1.regblock[16][10] ),
    .A1(\r1.regblock[17][10] ),
    .A2(\r1.regblock[18][10] ),
    .A3(\r1.regblock[19][10] ),
    .S0(net49),
    .S1(net42),
    .X(_00545_));
 sky130_fd_sc_hd__mux4_1 _14188_ (.A0(\r1.regblock[20][10] ),
    .A1(\r1.regblock[21][10] ),
    .A2(\r1.regblock[22][10] ),
    .A3(\r1.regblock[23][10] ),
    .S0(net49),
    .S1(net42),
    .X(_00546_));
 sky130_fd_sc_hd__mux4_1 _14189_ (.A0(\r1.regblock[24][10] ),
    .A1(\r1.regblock[25][10] ),
    .A2(\r1.regblock[26][10] ),
    .A3(\r1.regblock[27][10] ),
    .S0(net49),
    .S1(net42),
    .X(_00547_));
 sky130_fd_sc_hd__mux4_2 _14190_ (.A0(\r1.regblock[28][10] ),
    .A1(\r1.regblock[29][10] ),
    .A2(\r1.regblock[30][10] ),
    .A3(\r1.regblock[31][10] ),
    .S0(net49),
    .S1(net42),
    .X(_00548_));
 sky130_fd_sc_hd__mux4_2 _14191_ (.A0(_00545_),
    .A1(_00546_),
    .A2(_00547_),
    .A3(_00548_),
    .S0(net35),
    .S1(net33),
    .X(_00549_));
 sky130_fd_sc_hd__mux4_1 _14192_ (.A0(\r1.regblock[0][9] ),
    .A1(\r1.regblock[1][9] ),
    .A2(\r1.regblock[2][9] ),
    .A3(\r1.regblock[3][9] ),
    .S0(net48),
    .S1(net39),
    .X(_00527_));
 sky130_fd_sc_hd__mux4_2 _14193_ (.A0(\r1.regblock[4][9] ),
    .A1(\r1.regblock[5][9] ),
    .A2(\r1.regblock[6][9] ),
    .A3(\r1.regblock[7][9] ),
    .S0(net48),
    .S1(net39),
    .X(_00528_));
 sky130_fd_sc_hd__mux4_2 _14194_ (.A0(\r1.regblock[8][9] ),
    .A1(\r1.regblock[9][9] ),
    .A2(\r1.regblock[10][9] ),
    .A3(\r1.regblock[11][9] ),
    .S0(net48),
    .S1(net39),
    .X(_00529_));
 sky130_fd_sc_hd__mux4_1 _14195_ (.A0(\r1.regblock[12][9] ),
    .A1(\r1.regblock[13][9] ),
    .A2(\r1.regblock[14][9] ),
    .A3(\r1.regblock[15][9] ),
    .S0(net48),
    .S1(net39),
    .X(_00530_));
 sky130_fd_sc_hd__mux4_2 _14196_ (.A0(_00527_),
    .A1(_00528_),
    .A2(_00529_),
    .A3(_00530_),
    .S0(net35),
    .S1(net33),
    .X(_00531_));
 sky130_fd_sc_hd__mux4_1 _14197_ (.A0(\r1.regblock[16][9] ),
    .A1(\r1.regblock[17][9] ),
    .A2(\r1.regblock[18][9] ),
    .A3(\r1.regblock[19][9] ),
    .S0(net49),
    .S1(net42),
    .X(_00532_));
 sky130_fd_sc_hd__mux4_2 _14198_ (.A0(\r1.regblock[20][9] ),
    .A1(\r1.regblock[21][9] ),
    .A2(\r1.regblock[22][9] ),
    .A3(\r1.regblock[23][9] ),
    .S0(net49),
    .S1(net42),
    .X(_00533_));
 sky130_fd_sc_hd__mux4_1 _14199_ (.A0(\r1.regblock[24][9] ),
    .A1(\r1.regblock[25][9] ),
    .A2(\r1.regblock[26][9] ),
    .A3(\r1.regblock[27][9] ),
    .S0(net49),
    .S1(net42),
    .X(_00534_));
 sky130_fd_sc_hd__mux4_2 _14200_ (.A0(\r1.regblock[28][9] ),
    .A1(\r1.regblock[29][9] ),
    .A2(\r1.regblock[30][9] ),
    .A3(\r1.regblock[31][9] ),
    .S0(net49),
    .S1(net42),
    .X(_00535_));
 sky130_fd_sc_hd__mux4_2 _14201_ (.A0(_00532_),
    .A1(_00533_),
    .A2(_00534_),
    .A3(_00535_),
    .S0(net35),
    .S1(net33),
    .X(_00536_));
 sky130_fd_sc_hd__mux4_1 _14202_ (.A0(\r1.regblock[0][8] ),
    .A1(\r1.regblock[1][8] ),
    .A2(\r1.regblock[2][8] ),
    .A3(\r1.regblock[3][8] ),
    .S0(net48),
    .S1(net39),
    .X(_00514_));
 sky130_fd_sc_hd__mux4_2 _14203_ (.A0(\r1.regblock[4][8] ),
    .A1(\r1.regblock[5][8] ),
    .A2(\r1.regblock[6][8] ),
    .A3(\r1.regblock[7][8] ),
    .S0(net48),
    .S1(net39),
    .X(_00515_));
 sky130_fd_sc_hd__mux4_2 _14204_ (.A0(\r1.regblock[8][8] ),
    .A1(\r1.regblock[9][8] ),
    .A2(\r1.regblock[10][8] ),
    .A3(\r1.regblock[11][8] ),
    .S0(net48),
    .S1(net39),
    .X(_00516_));
 sky130_fd_sc_hd__mux4_2 _14205_ (.A0(\r1.regblock[12][8] ),
    .A1(\r1.regblock[13][8] ),
    .A2(\r1.regblock[14][8] ),
    .A3(\r1.regblock[15][8] ),
    .S0(net48),
    .S1(net39),
    .X(_00517_));
 sky130_fd_sc_hd__mux4_2 _14206_ (.A0(_00514_),
    .A1(_00515_),
    .A2(_00516_),
    .A3(_00517_),
    .S0(net35),
    .S1(net33),
    .X(_00518_));
 sky130_fd_sc_hd__mux4_1 _14207_ (.A0(\r1.regblock[16][8] ),
    .A1(\r1.regblock[17][8] ),
    .A2(\r1.regblock[18][8] ),
    .A3(\r1.regblock[19][8] ),
    .S0(net49),
    .S1(net42),
    .X(_00519_));
 sky130_fd_sc_hd__mux4_2 _14208_ (.A0(\r1.regblock[20][8] ),
    .A1(\r1.regblock[21][8] ),
    .A2(\r1.regblock[22][8] ),
    .A3(\r1.regblock[23][8] ),
    .S0(net49),
    .S1(net42),
    .X(_00520_));
 sky130_fd_sc_hd__mux4_1 _14209_ (.A0(\r1.regblock[24][8] ),
    .A1(\r1.regblock[25][8] ),
    .A2(\r1.regblock[26][8] ),
    .A3(\r1.regblock[27][8] ),
    .S0(net49),
    .S1(net42),
    .X(_00521_));
 sky130_fd_sc_hd__mux4_2 _14210_ (.A0(\r1.regblock[28][8] ),
    .A1(\r1.regblock[29][8] ),
    .A2(\r1.regblock[30][8] ),
    .A3(\r1.regblock[31][8] ),
    .S0(net49),
    .S1(net42),
    .X(_00522_));
 sky130_fd_sc_hd__mux4_2 _14211_ (.A0(_00519_),
    .A1(_00520_),
    .A2(_00521_),
    .A3(_00522_),
    .S0(net35),
    .S1(net33),
    .X(_00523_));
 sky130_fd_sc_hd__mux4_2 _14212_ (.A0(\r1.regblock[0][7] ),
    .A1(\r1.regblock[1][7] ),
    .A2(\r1.regblock[2][7] ),
    .A3(\r1.regblock[3][7] ),
    .S0(net48),
    .S1(net39),
    .X(_00501_));
 sky130_fd_sc_hd__mux4_2 _14213_ (.A0(\r1.regblock[4][7] ),
    .A1(\r1.regblock[5][7] ),
    .A2(\r1.regblock[6][7] ),
    .A3(\r1.regblock[7][7] ),
    .S0(net48),
    .S1(net39),
    .X(_00502_));
 sky130_fd_sc_hd__mux4_1 _14214_ (.A0(\r1.regblock[8][7] ),
    .A1(\r1.regblock[9][7] ),
    .A2(\r1.regblock[10][7] ),
    .A3(\r1.regblock[11][7] ),
    .S0(net48),
    .S1(net39),
    .X(_00503_));
 sky130_fd_sc_hd__mux4_1 _14215_ (.A0(\r1.regblock[12][7] ),
    .A1(\r1.regblock[13][7] ),
    .A2(\r1.regblock[14][7] ),
    .A3(\r1.regblock[15][7] ),
    .S0(net48),
    .S1(net39),
    .X(_00504_));
 sky130_fd_sc_hd__mux4_2 _14216_ (.A0(_00501_),
    .A1(_00502_),
    .A2(_00503_),
    .A3(_00504_),
    .S0(net35),
    .S1(net33),
    .X(_00505_));
 sky130_fd_sc_hd__mux4_1 _14217_ (.A0(\r1.regblock[16][7] ),
    .A1(\r1.regblock[17][7] ),
    .A2(\r1.regblock[18][7] ),
    .A3(\r1.regblock[19][7] ),
    .S0(net49),
    .S1(net40),
    .X(_00506_));
 sky130_fd_sc_hd__mux4_2 _14218_ (.A0(\r1.regblock[20][7] ),
    .A1(\r1.regblock[21][7] ),
    .A2(\r1.regblock[22][7] ),
    .A3(\r1.regblock[23][7] ),
    .S0(net49),
    .S1(net40),
    .X(_00507_));
 sky130_fd_sc_hd__mux4_2 _14219_ (.A0(\r1.regblock[24][7] ),
    .A1(\r1.regblock[25][7] ),
    .A2(\r1.regblock[26][7] ),
    .A3(\r1.regblock[27][7] ),
    .S0(net48),
    .S1(net39),
    .X(_00508_));
 sky130_fd_sc_hd__mux4_2 _14220_ (.A0(\r1.regblock[28][7] ),
    .A1(\r1.regblock[29][7] ),
    .A2(\r1.regblock[30][7] ),
    .A3(\r1.regblock[31][7] ),
    .S0(net48),
    .S1(net39),
    .X(_00509_));
 sky130_fd_sc_hd__mux4_1 _14221_ (.A0(_00506_),
    .A1(_00507_),
    .A2(_00508_),
    .A3(_00509_),
    .S0(net35),
    .S1(net33),
    .X(_00510_));
 sky130_fd_sc_hd__mux4_1 _14222_ (.A0(\r1.regblock[0][6] ),
    .A1(\r1.regblock[1][6] ),
    .A2(\r1.regblock[2][6] ),
    .A3(\r1.regblock[3][6] ),
    .S0(net47),
    .S1(net39),
    .X(_00488_));
 sky130_fd_sc_hd__mux4_2 _14223_ (.A0(\r1.regblock[4][6] ),
    .A1(\r1.regblock[5][6] ),
    .A2(\r1.regblock[6][6] ),
    .A3(\r1.regblock[7][6] ),
    .S0(net47),
    .S1(net39),
    .X(_00489_));
 sky130_fd_sc_hd__mux4_2 _14224_ (.A0(\r1.regblock[8][6] ),
    .A1(\r1.regblock[9][6] ),
    .A2(\r1.regblock[10][6] ),
    .A3(\r1.regblock[11][6] ),
    .S0(net48),
    .S1(net39),
    .X(_00490_));
 sky130_fd_sc_hd__mux4_1 _14225_ (.A0(\r1.regblock[12][6] ),
    .A1(\r1.regblock[13][6] ),
    .A2(\r1.regblock[14][6] ),
    .A3(\r1.regblock[15][6] ),
    .S0(net47),
    .S1(net39),
    .X(_00491_));
 sky130_fd_sc_hd__mux4_2 _14226_ (.A0(_00488_),
    .A1(_00489_),
    .A2(_00490_),
    .A3(_00491_),
    .S0(net35),
    .S1(net33),
    .X(_00492_));
 sky130_fd_sc_hd__mux4_1 _14227_ (.A0(\r1.regblock[16][6] ),
    .A1(\r1.regblock[17][6] ),
    .A2(\r1.regblock[18][6] ),
    .A3(\r1.regblock[19][6] ),
    .S0(net49),
    .S1(net40),
    .X(_00493_));
 sky130_fd_sc_hd__mux4_2 _14228_ (.A0(\r1.regblock[20][6] ),
    .A1(\r1.regblock[21][6] ),
    .A2(\r1.regblock[22][6] ),
    .A3(\r1.regblock[23][6] ),
    .S0(net46),
    .S1(net41),
    .X(_00494_));
 sky130_fd_sc_hd__mux4_2 _14229_ (.A0(\r1.regblock[24][6] ),
    .A1(\r1.regblock[25][6] ),
    .A2(\r1.regblock[26][6] ),
    .A3(\r1.regblock[27][6] ),
    .S0(net48),
    .S1(net39),
    .X(_00495_));
 sky130_fd_sc_hd__mux4_1 _14230_ (.A0(\r1.regblock[28][6] ),
    .A1(\r1.regblock[29][6] ),
    .A2(\r1.regblock[30][6] ),
    .A3(\r1.regblock[31][6] ),
    .S0(net49),
    .S1(net40),
    .X(_00496_));
 sky130_fd_sc_hd__mux4_1 _14231_ (.A0(_00493_),
    .A1(_00494_),
    .A2(_00495_),
    .A3(_00496_),
    .S0(net35),
    .S1(net33),
    .X(_00497_));
 sky130_fd_sc_hd__mux4_2 _14232_ (.A0(\r1.regblock[0][5] ),
    .A1(\r1.regblock[1][5] ),
    .A2(\r1.regblock[2][5] ),
    .A3(\r1.regblock[3][5] ),
    .S0(net47),
    .S1(net39),
    .X(_00475_));
 sky130_fd_sc_hd__mux4_2 _14233_ (.A0(\r1.regblock[4][5] ),
    .A1(\r1.regblock[5][5] ),
    .A2(\r1.regblock[6][5] ),
    .A3(\r1.regblock[7][5] ),
    .S0(net47),
    .S1(net39),
    .X(_00476_));
 sky130_fd_sc_hd__mux4_1 _14234_ (.A0(\r1.regblock[8][5] ),
    .A1(\r1.regblock[9][5] ),
    .A2(\r1.regblock[10][5] ),
    .A3(\r1.regblock[11][5] ),
    .S0(net47),
    .S1(net39),
    .X(_00477_));
 sky130_fd_sc_hd__mux4_1 _14235_ (.A0(\r1.regblock[12][5] ),
    .A1(\r1.regblock[13][5] ),
    .A2(\r1.regblock[14][5] ),
    .A3(\r1.regblock[15][5] ),
    .S0(net47),
    .S1(net39),
    .X(_00478_));
 sky130_fd_sc_hd__mux4_2 _14236_ (.A0(_00475_),
    .A1(_00476_),
    .A2(_00477_),
    .A3(_00478_),
    .S0(net35),
    .S1(net33),
    .X(_00479_));
 sky130_fd_sc_hd__mux4_1 _14237_ (.A0(\r1.regblock[16][5] ),
    .A1(\r1.regblock[17][5] ),
    .A2(\r1.regblock[18][5] ),
    .A3(\r1.regblock[19][5] ),
    .S0(net49),
    .S1(net40),
    .X(_00480_));
 sky130_fd_sc_hd__mux4_2 _14238_ (.A0(\r1.regblock[20][5] ),
    .A1(\r1.regblock[21][5] ),
    .A2(\r1.regblock[22][5] ),
    .A3(\r1.regblock[23][5] ),
    .S0(net46),
    .S1(net41),
    .X(_00481_));
 sky130_fd_sc_hd__mux4_2 _14239_ (.A0(\r1.regblock[24][5] ),
    .A1(\r1.regblock[25][5] ),
    .A2(\r1.regblock[26][5] ),
    .A3(\r1.regblock[27][5] ),
    .S0(net48),
    .S1(net39),
    .X(_00482_));
 sky130_fd_sc_hd__mux4_2 _14240_ (.A0(\r1.regblock[28][5] ),
    .A1(\r1.regblock[29][5] ),
    .A2(\r1.regblock[30][5] ),
    .A3(\r1.regblock[31][5] ),
    .S0(net49),
    .S1(net40),
    .X(_00483_));
 sky130_fd_sc_hd__mux4_1 _14241_ (.A0(_00480_),
    .A1(_00481_),
    .A2(_00482_),
    .A3(_00483_),
    .S0(net35),
    .S1(net32),
    .X(_00484_));
 sky130_fd_sc_hd__mux4_2 _14242_ (.A0(\r1.regblock[0][4] ),
    .A1(\r1.regblock[1][4] ),
    .A2(\r1.regblock[2][4] ),
    .A3(\r1.regblock[3][4] ),
    .S0(net47),
    .S1(net39),
    .X(_00462_));
 sky130_fd_sc_hd__mux4_2 _14243_ (.A0(\r1.regblock[4][4] ),
    .A1(\r1.regblock[5][4] ),
    .A2(\r1.regblock[6][4] ),
    .A3(\r1.regblock[7][4] ),
    .S0(net47),
    .S1(net39),
    .X(_00463_));
 sky130_fd_sc_hd__mux4_1 _14244_ (.A0(\r1.regblock[8][4] ),
    .A1(\r1.regblock[9][4] ),
    .A2(\r1.regblock[10][4] ),
    .A3(\r1.regblock[11][4] ),
    .S0(net47),
    .S1(net39),
    .X(_00464_));
 sky130_fd_sc_hd__mux4_1 _14245_ (.A0(\r1.regblock[12][4] ),
    .A1(\r1.regblock[13][4] ),
    .A2(\r1.regblock[14][4] ),
    .A3(\r1.regblock[15][4] ),
    .S0(net47),
    .S1(net39),
    .X(_00465_));
 sky130_fd_sc_hd__mux4_2 _14246_ (.A0(_00462_),
    .A1(_00463_),
    .A2(_00464_),
    .A3(_00465_),
    .S0(net35),
    .S1(net33),
    .X(_00466_));
 sky130_fd_sc_hd__mux4_1 _14247_ (.A0(\r1.regblock[16][4] ),
    .A1(\r1.regblock[17][4] ),
    .A2(\r1.regblock[18][4] ),
    .A3(\r1.regblock[19][4] ),
    .S0(net49),
    .S1(net40),
    .X(_00467_));
 sky130_fd_sc_hd__mux4_2 _14248_ (.A0(\r1.regblock[20][4] ),
    .A1(\r1.regblock[21][4] ),
    .A2(\r1.regblock[22][4] ),
    .A3(\r1.regblock[23][4] ),
    .S0(net49),
    .S1(net40),
    .X(_00468_));
 sky130_fd_sc_hd__mux4_1 _14249_ (.A0(\r1.regblock[24][4] ),
    .A1(\r1.regblock[25][4] ),
    .A2(\r1.regblock[26][4] ),
    .A3(\r1.regblock[27][4] ),
    .S0(net49),
    .S1(net40),
    .X(_00469_));
 sky130_fd_sc_hd__mux4_2 _14250_ (.A0(\r1.regblock[28][4] ),
    .A1(\r1.regblock[29][4] ),
    .A2(\r1.regblock[30][4] ),
    .A3(\r1.regblock[31][4] ),
    .S0(net50),
    .S1(net40),
    .X(_00470_));
 sky130_fd_sc_hd__mux4_1 _14251_ (.A0(_00467_),
    .A1(_00468_),
    .A2(_00469_),
    .A3(_00470_),
    .S0(net34),
    .S1(net32),
    .X(_00471_));
 sky130_fd_sc_hd__mux4_2 _14252_ (.A0(\r1.regblock[0][3] ),
    .A1(\r1.regblock[1][3] ),
    .A2(\r1.regblock[2][3] ),
    .A3(\r1.regblock[3][3] ),
    .S0(net47),
    .S1(net39),
    .X(_00449_));
 sky130_fd_sc_hd__mux4_2 _14253_ (.A0(\r1.regblock[4][3] ),
    .A1(\r1.regblock[5][3] ),
    .A2(\r1.regblock[6][3] ),
    .A3(\r1.regblock[7][3] ),
    .S0(net47),
    .S1(net39),
    .X(_00450_));
 sky130_fd_sc_hd__mux4_1 _14254_ (.A0(\r1.regblock[8][3] ),
    .A1(\r1.regblock[9][3] ),
    .A2(\r1.regblock[10][3] ),
    .A3(\r1.regblock[11][3] ),
    .S0(net47),
    .S1(net39),
    .X(_00451_));
 sky130_fd_sc_hd__mux4_1 _14255_ (.A0(\r1.regblock[12][3] ),
    .A1(\r1.regblock[13][3] ),
    .A2(\r1.regblock[14][3] ),
    .A3(\r1.regblock[15][3] ),
    .S0(net47),
    .S1(net39),
    .X(_00452_));
 sky130_fd_sc_hd__mux4_2 _14256_ (.A0(_00449_),
    .A1(_00450_),
    .A2(_00451_),
    .A3(_00452_),
    .S0(net35),
    .S1(net33),
    .X(_00453_));
 sky130_fd_sc_hd__mux4_1 _14257_ (.A0(\r1.regblock[16][3] ),
    .A1(\r1.regblock[17][3] ),
    .A2(\r1.regblock[18][3] ),
    .A3(\r1.regblock[19][3] ),
    .S0(net50),
    .S1(net40),
    .X(_00454_));
 sky130_fd_sc_hd__mux4_2 _14258_ (.A0(\r1.regblock[20][3] ),
    .A1(\r1.regblock[21][3] ),
    .A2(\r1.regblock[22][3] ),
    .A3(\r1.regblock[23][3] ),
    .S0(net49),
    .S1(net40),
    .X(_00455_));
 sky130_fd_sc_hd__mux4_1 _14259_ (.A0(\r1.regblock[24][3] ),
    .A1(\r1.regblock[25][3] ),
    .A2(\r1.regblock[26][3] ),
    .A3(\r1.regblock[27][3] ),
    .S0(net50),
    .S1(net40),
    .X(_00456_));
 sky130_fd_sc_hd__mux4_2 _14260_ (.A0(\r1.regblock[28][3] ),
    .A1(\r1.regblock[29][3] ),
    .A2(\r1.regblock[30][3] ),
    .A3(\r1.regblock[31][3] ),
    .S0(net50),
    .S1(net40),
    .X(_00457_));
 sky130_fd_sc_hd__mux4_1 _14261_ (.A0(_00454_),
    .A1(_00455_),
    .A2(_00456_),
    .A3(_00457_),
    .S0(net34),
    .S1(net32),
    .X(_00458_));
 sky130_fd_sc_hd__mux4_1 _14262_ (.A0(\r1.regblock[0][2] ),
    .A1(\r1.regblock[1][2] ),
    .A2(\r1.regblock[2][2] ),
    .A3(\r1.regblock[3][2] ),
    .S0(net47),
    .S1(net39),
    .X(_00436_));
 sky130_fd_sc_hd__mux4_2 _14263_ (.A0(\r1.regblock[4][2] ),
    .A1(\r1.regblock[5][2] ),
    .A2(\r1.regblock[6][2] ),
    .A3(\r1.regblock[7][2] ),
    .S0(net47),
    .S1(net39),
    .X(_00437_));
 sky130_fd_sc_hd__mux4_1 _14264_ (.A0(\r1.regblock[8][2] ),
    .A1(\r1.regblock[9][2] ),
    .A2(\r1.regblock[10][2] ),
    .A3(\r1.regblock[11][2] ),
    .S0(net47),
    .S1(net39),
    .X(_00438_));
 sky130_fd_sc_hd__mux4_2 _14265_ (.A0(\r1.regblock[12][2] ),
    .A1(\r1.regblock[13][2] ),
    .A2(\r1.regblock[14][2] ),
    .A3(\r1.regblock[15][2] ),
    .S0(net47),
    .S1(net39),
    .X(_00439_));
 sky130_fd_sc_hd__mux4_2 _14266_ (.A0(_00436_),
    .A1(_00437_),
    .A2(_00438_),
    .A3(_00439_),
    .S0(net35),
    .S1(net33),
    .X(_00440_));
 sky130_fd_sc_hd__mux4_1 _14267_ (.A0(\r1.regblock[16][2] ),
    .A1(\r1.regblock[17][2] ),
    .A2(\r1.regblock[18][2] ),
    .A3(\r1.regblock[19][2] ),
    .S0(net50),
    .S1(net40),
    .X(_00441_));
 sky130_fd_sc_hd__mux4_2 _14268_ (.A0(\r1.regblock[20][2] ),
    .A1(\r1.regblock[21][2] ),
    .A2(\r1.regblock[22][2] ),
    .A3(\r1.regblock[23][2] ),
    .S0(net49),
    .S1(net40),
    .X(_00442_));
 sky130_fd_sc_hd__mux4_1 _14269_ (.A0(\r1.regblock[24][2] ),
    .A1(\r1.regblock[25][2] ),
    .A2(\r1.regblock[26][2] ),
    .A3(\r1.regblock[27][2] ),
    .S0(net50),
    .S1(net40),
    .X(_00443_));
 sky130_fd_sc_hd__mux4_2 _14270_ (.A0(\r1.regblock[28][2] ),
    .A1(\r1.regblock[29][2] ),
    .A2(\r1.regblock[30][2] ),
    .A3(\r1.regblock[31][2] ),
    .S0(net50),
    .S1(net40),
    .X(_00444_));
 sky130_fd_sc_hd__mux4_1 _14271_ (.A0(_00441_),
    .A1(_00442_),
    .A2(_00443_),
    .A3(_00444_),
    .S0(net34),
    .S1(net32),
    .X(_00445_));
 sky130_fd_sc_hd__mux4_2 _14272_ (.A0(\r1.regblock[0][1] ),
    .A1(\r1.regblock[1][1] ),
    .A2(\r1.regblock[2][1] ),
    .A3(\r1.regblock[3][1] ),
    .S0(net50),
    .S1(net40),
    .X(_00423_));
 sky130_fd_sc_hd__mux4_2 _14273_ (.A0(\r1.regblock[4][1] ),
    .A1(\r1.regblock[5][1] ),
    .A2(\r1.regblock[6][1] ),
    .A3(\r1.regblock[7][1] ),
    .S0(net43),
    .S1(net38),
    .X(_00424_));
 sky130_fd_sc_hd__mux4_1 _14274_ (.A0(\r1.regblock[8][1] ),
    .A1(\r1.regblock[9][1] ),
    .A2(\r1.regblock[10][1] ),
    .A3(\r1.regblock[11][1] ),
    .S0(net50),
    .S1(net40),
    .X(_00425_));
 sky130_fd_sc_hd__mux4_1 _14275_ (.A0(\r1.regblock[12][1] ),
    .A1(\r1.regblock[13][1] ),
    .A2(\r1.regblock[14][1] ),
    .A3(\r1.regblock[15][1] ),
    .S0(net50),
    .S1(net40),
    .X(_00426_));
 sky130_fd_sc_hd__mux4_2 _14276_ (.A0(_00423_),
    .A1(_00424_),
    .A2(_00425_),
    .A3(_00426_),
    .S0(net34),
    .S1(net32),
    .X(_00427_));
 sky130_fd_sc_hd__mux4_2 _14277_ (.A0(\r1.regblock[16][1] ),
    .A1(\r1.regblock[17][1] ),
    .A2(\r1.regblock[18][1] ),
    .A3(\r1.regblock[19][1] ),
    .S0(net50),
    .S1(net40),
    .X(_00428_));
 sky130_fd_sc_hd__mux4_2 _14278_ (.A0(\r1.regblock[20][1] ),
    .A1(\r1.regblock[21][1] ),
    .A2(\r1.regblock[22][1] ),
    .A3(\r1.regblock[23][1] ),
    .S0(net50),
    .S1(net40),
    .X(_00429_));
 sky130_fd_sc_hd__mux4_1 _14279_ (.A0(\r1.regblock[24][1] ),
    .A1(\r1.regblock[25][1] ),
    .A2(\r1.regblock[26][1] ),
    .A3(\r1.regblock[27][1] ),
    .S0(net50),
    .S1(net40),
    .X(_00430_));
 sky130_fd_sc_hd__mux4_2 _14280_ (.A0(\r1.regblock[28][1] ),
    .A1(\r1.regblock[29][1] ),
    .A2(\r1.regblock[30][1] ),
    .A3(\r1.regblock[31][1] ),
    .S0(net50),
    .S1(net40),
    .X(_00431_));
 sky130_fd_sc_hd__mux4_1 _14281_ (.A0(_00428_),
    .A1(_00429_),
    .A2(_00430_),
    .A3(_00431_),
    .S0(\c1.instruction1[22] ),
    .S1(\c1.instruction1[23] ),
    .X(_00432_));
 sky130_fd_sc_hd__mux4_1 _14282_ (.A0(\r1.regblock[0][0] ),
    .A1(\r1.regblock[1][0] ),
    .A2(\r1.regblock[2][0] ),
    .A3(\r1.regblock[3][0] ),
    .S0(net50),
    .S1(net40),
    .X(_00409_));
 sky130_fd_sc_hd__mux4_2 _14283_ (.A0(\r1.regblock[4][0] ),
    .A1(\r1.regblock[5][0] ),
    .A2(\r1.regblock[6][0] ),
    .A3(\r1.regblock[7][0] ),
    .S0(net43),
    .S1(net38),
    .X(_00410_));
 sky130_fd_sc_hd__mux4_1 _14284_ (.A0(\r1.regblock[8][0] ),
    .A1(\r1.regblock[9][0] ),
    .A2(\r1.regblock[10][0] ),
    .A3(\r1.regblock[11][0] ),
    .S0(net50),
    .S1(net38),
    .X(_00411_));
 sky130_fd_sc_hd__mux4_1 _14285_ (.A0(\r1.regblock[12][0] ),
    .A1(\r1.regblock[13][0] ),
    .A2(\r1.regblock[14][0] ),
    .A3(\r1.regblock[15][0] ),
    .S0(net50),
    .S1(net40),
    .X(_00412_));
 sky130_fd_sc_hd__mux4_2 _14286_ (.A0(_00409_),
    .A1(_00410_),
    .A2(_00411_),
    .A3(_00412_),
    .S0(net34),
    .S1(net32),
    .X(_00413_));
 sky130_fd_sc_hd__mux4_1 _14287_ (.A0(\r1.regblock[16][0] ),
    .A1(\r1.regblock[17][0] ),
    .A2(\r1.regblock[18][0] ),
    .A3(\r1.regblock[19][0] ),
    .S0(net50),
    .S1(net40),
    .X(_00414_));
 sky130_fd_sc_hd__mux4_1 _14288_ (.A0(\r1.regblock[20][0] ),
    .A1(\r1.regblock[21][0] ),
    .A2(\r1.regblock[22][0] ),
    .A3(\r1.regblock[23][0] ),
    .S0(net50),
    .S1(net40),
    .X(_00415_));
 sky130_fd_sc_hd__mux4_1 _14289_ (.A0(\r1.regblock[24][0] ),
    .A1(\r1.regblock[25][0] ),
    .A2(\r1.regblock[26][0] ),
    .A3(\r1.regblock[27][0] ),
    .S0(net50),
    .S1(net40),
    .X(_00416_));
 sky130_fd_sc_hd__mux4_2 _14290_ (.A0(\r1.regblock[28][0] ),
    .A1(\r1.regblock[29][0] ),
    .A2(\r1.regblock[30][0] ),
    .A3(\r1.regblock[31][0] ),
    .S0(net50),
    .S1(net40),
    .X(_00417_));
 sky130_fd_sc_hd__mux4_1 _14291_ (.A0(_00414_),
    .A1(_00415_),
    .A2(_00416_),
    .A3(_00417_),
    .S0(\c1.instruction1[22] ),
    .S1(\c1.instruction1[23] ),
    .X(_00418_));
 sky130_fd_sc_hd__dfxtp_1 _14292_ (.D(\c1.instruction3[0] ),
    .Q(\w1.instruction[0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _14293_ (.D(\c1.instruction3[1] ),
    .Q(\w1.instruction[1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _14294_ (.D(\c1.instruction3[2] ),
    .Q(\w1.instruction[2] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _14295_ (.D(\c1.instruction3[3] ),
    .Q(\w1.instruction[3] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _14296_ (.D(\c1.instruction3[4] ),
    .Q(\w1.instruction[4] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _14297_ (.D(\c1.instruction3[5] ),
    .Q(\w1.instruction[5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _14298_ (.D(\c1.instruction3[6] ),
    .Q(\w1.instruction[6] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _14299_ (.D(\c1.instruction3[7] ),
    .Q(\r1.waddr[0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _14300_ (.D(\c1.instruction3[8] ),
    .Q(\r1.waddr[1] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _14301_ (.D(\c1.instruction3[9] ),
    .Q(\r1.waddr[2] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _14302_ (.D(\c1.instruction3[10] ),
    .Q(\r1.waddr[3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _14303_ (.D(\c1.instruction3[11] ),
    .Q(\r1.waddr[4] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _14304_ (.D(\wbmemout[0] ),
    .Q(\r1.wdata[0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 _14305_ (.D(\wbmemout[1] ),
    .Q(\r1.wdata[1] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _14306_ (.D(\wbmemout[2] ),
    .Q(\r1.wdata[2] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _14307_ (.D(\wbmemout[3] ),
    .Q(\r1.wdata[3] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_2 _14308_ (.D(\wbmemout[4] ),
    .Q(\r1.wdata[4] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 _14309_ (.D(\wbmemout[5] ),
    .Q(\r1.wdata[5] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _14310_ (.D(\wbmemout[6] ),
    .Q(\r1.wdata[6] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _14311_ (.D(\wbmemout[7] ),
    .Q(\r1.wdata[7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _14312_ (.D(\wbmemout[8] ),
    .Q(\r1.wdata[8] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _14313_ (.D(\wbmemout[9] ),
    .Q(\r1.wdata[9] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _14314_ (.D(\wbmemout[10] ),
    .Q(\r1.wdata[10] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _14315_ (.D(\wbmemout[11] ),
    .Q(\r1.wdata[11] ),
    .CLK(clknet_2_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _14316_ (.D(\wbmemout[12] ),
    .Q(\r1.wdata[12] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 _14317_ (.D(\wbmemout[13] ),
    .Q(\r1.wdata[13] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 _14318_ (.D(\wbmemout[14] ),
    .Q(\r1.wdata[14] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 _14319_ (.D(\wbmemout[15] ),
    .Q(\r1.wdata[15] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _14320_ (.D(\wbmemout[16] ),
    .Q(\r1.wdata[16] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _14321_ (.D(\wbmemout[17] ),
    .Q(\r1.wdata[17] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _14322_ (.D(\wbmemout[18] ),
    .Q(\r1.wdata[18] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 _14323_ (.D(\wbmemout[19] ),
    .Q(\r1.wdata[19] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _14324_ (.D(\wbmemout[20] ),
    .Q(\r1.wdata[20] ),
    .CLK(clknet_opt_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _14325_ (.D(\wbmemout[21] ),
    .Q(\r1.wdata[21] ),
    .CLK(clknet_2_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _14326_ (.D(\wbmemout[22] ),
    .Q(\r1.wdata[22] ),
    .CLK(clknet_2_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _14327_ (.D(\wbmemout[23] ),
    .Q(\r1.wdata[23] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 _14328_ (.D(\wbmemout[24] ),
    .Q(\r1.wdata[24] ),
    .CLK(clknet_2_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _14329_ (.D(\wbmemout[25] ),
    .Q(\r1.wdata[25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _14330_ (.D(\wbmemout[26] ),
    .Q(\r1.wdata[26] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _14331_ (.D(\wbmemout[27] ),
    .Q(\r1.wdata[27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 _14332_ (.D(\wbmemout[28] ),
    .Q(\r1.wdata[28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _14333_ (.D(\wbmemout[29] ),
    .Q(\r1.wdata[29] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 _14334_ (.D(\wbmemout[30] ),
    .Q(\r1.wdata[30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _14335_ (.D(\wbmemout[31] ),
    .Q(\r1.wdata[31] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_4 _14336_ (.D(\c1.dep_place[0] ),
    .Q(\DEP_PLACE[0] ),
    .CLK(_01369_));
 sky130_fd_sc_hd__dfxtp_4 _14337_ (.D(\c1.dep_place[1] ),
    .Q(\DEP_PLACE[1] ),
    .CLK(_01370_));
 sky130_fd_sc_hd__dfxtp_4 _14338_ (.D(\c1.dep_place[2] ),
    .Q(\DEP_PLACE[2] ),
    .CLK(_01371_));
 sky130_fd_sc_hd__dfxtp_1 _14339_ (.D(pc[0]),
    .Q(\e1.pc[0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _14340_ (.D(pc[1]),
    .Q(\e1.pc[1] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _14341_ (.D(pc[2]),
    .Q(\e1.pc[2] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 _14342_ (.D(pc[3]),
    .Q(\e1.pc[3] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _14343_ (.D(pc[4]),
    .Q(\e1.pc[4] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _14344_ (.D(pc[5]),
    .Q(\e1.pc[5] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _14345_ (.D(pc[6]),
    .Q(\e1.pc[6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _14346_ (.D(pc[7]),
    .Q(\e1.pc[7] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _14347_ (.D(pc[8]),
    .Q(\e1.pc[8] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _14348_ (.D(pc[9]),
    .Q(\e1.pc[9] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _14349_ (.D(pc[10]),
    .Q(\e1.pc[10] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _14350_ (.D(pc[11]),
    .Q(\e1.pc[11] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _14351_ (.D(pc[12]),
    .Q(\e1.pc[12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _14352_ (.D(pc[13]),
    .Q(\e1.pc[13] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _14353_ (.D(pc[14]),
    .Q(\e1.pc[14] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _14354_ (.D(pc[15]),
    .Q(\e1.pc[15] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _14355_ (.D(pc[16]),
    .Q(\e1.pc[16] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _14356_ (.D(pc[17]),
    .Q(\e1.pc[17] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _14357_ (.D(pc[18]),
    .Q(\e1.pc[18] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _14358_ (.D(pc[19]),
    .Q(\e1.pc[19] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _14359_ (.D(pc[20]),
    .Q(\e1.pc[20] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _14360_ (.D(pc[21]),
    .Q(\e1.pc[21] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _14361_ (.D(pc[22]),
    .Q(\e1.pc[22] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _14362_ (.D(pc[23]),
    .Q(\e1.pc[23] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _14363_ (.D(pc[24]),
    .Q(\e1.pc[24] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 _14364_ (.D(pc[25]),
    .Q(\e1.pc[25] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 _14365_ (.D(pc[26]),
    .Q(\e1.pc[26] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 _14366_ (.D(pc[27]),
    .Q(\e1.pc[27] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _14367_ (.D(pc[28]),
    .Q(\e1.pc[28] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _14368_ (.D(pc[29]),
    .Q(\e1.pc[29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _14369_ (.D(pc[30]),
    .Q(\e1.pc[30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _14370_ (.D(pc[31]),
    .Q(\e1.pc[31] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_4 _14371_ (.D(instruction[0]),
    .Q(\c1.instruction1[0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _14372_ (.D(instruction[1]),
    .Q(\c1.instruction1[1] ),
    .CLK(clknet_opt_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _14373_ (.D(instruction[2]),
    .Q(\c1.instruction1[2] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _14374_ (.D(instruction[3]),
    .Q(\c1.instruction1[3] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 _14375_ (.D(instruction[4]),
    .Q(\c1.instruction1[4] ),
    .CLK(clknet_opt_1_clk));
 sky130_fd_sc_hd__dfxtp_2 _14376_ (.D(instruction[5]),
    .Q(\c1.instruction1[5] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 _14377_ (.D(instruction[6]),
    .Q(\c1.instruction1[6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 _14378_ (.D(instruction[7]),
    .Q(\c1.instruction1[7] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_2 _14379_ (.D(instruction[8]),
    .Q(\c1.instruction1[8] ),
    .CLK(clknet_opt_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _14380_ (.D(instruction[9]),
    .Q(\c1.instruction1[9] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_2 _14381_ (.D(instruction[10]),
    .Q(\c1.instruction1[10] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_2 _14382_ (.D(instruction[11]),
    .Q(\c1.instruction1[11] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_4 _14383_ (.D(instruction[12]),
    .Q(\c1.instruction1[12] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _14384_ (.D(instruction[13]),
    .Q(\c1.instruction1[13] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_2 _14385_ (.D(instruction[14]),
    .Q(\c1.instruction1[14] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_4 _14386_ (.D(instruction[19]),
    .Q(\c1.instruction1[19] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_4 _14387_ (.D(instruction[24]),
    .Q(\c1.instruction1[24] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_4 _14388_ (.D(instruction[25]),
    .Q(\c1.instruction1[25] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_2 _14389_ (.D(instruction[26]),
    .Q(\c1.instruction1[26] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _14390_ (.D(instruction[27]),
    .Q(\c1.instruction1[27] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_2 _14391_ (.D(instruction[28]),
    .Q(\c1.instruction1[28] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_2 _14392_ (.D(instruction[29]),
    .Q(\c1.instruction1[29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_2 _14393_ (.D(instruction[30]),
    .Q(\c1.instruction1[30] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_4 _14394_ (.D(instruction[31]),
    .Q(\c1.instruction1[31] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_4 _14395_ (.D(instruction[20]),
    .Q(\c1.instruction1[20] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_4 _14396_ (.D(instruction[21]),
    .Q(\c1.instruction1[21] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 _14397_ (.D(instruction[22]),
    .Q(\c1.instruction1[22] ),
    .CLK(clknet_2_2_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _14398_ (.D(instruction[23]),
    .Q(\c1.instruction1[23] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_4 _14399_ (.D(instruction[15]),
    .Q(\c1.instruction1[15] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_4 _14400_ (.D(instruction[16]),
    .Q(\c1.instruction1[16] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_4 _14401_ (.D(instruction[17]),
    .Q(\c1.instruction1[17] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_4 _14402_ (.D(instruction[18]),
    .Q(\c1.instruction1[18] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _14403_ (.D(_02397_),
    .Q(\r1.regblock[23][0] ),
    .CLK(_01372_));
 sky130_fd_sc_hd__dfxtp_1 _14404_ (.D(_02398_),
    .Q(\r1.regblock[23][1] ),
    .CLK(_01373_));
 sky130_fd_sc_hd__dfxtp_1 _14405_ (.D(_02399_),
    .Q(\r1.regblock[23][2] ),
    .CLK(_01374_));
 sky130_fd_sc_hd__dfxtp_1 _14406_ (.D(_02400_),
    .Q(\r1.regblock[23][3] ),
    .CLK(_01375_));
 sky130_fd_sc_hd__dfxtp_1 _14407_ (.D(_02401_),
    .Q(\r1.regblock[23][4] ),
    .CLK(_01376_));
 sky130_fd_sc_hd__dfxtp_1 _14408_ (.D(_02402_),
    .Q(\r1.regblock[23][5] ),
    .CLK(_01377_));
 sky130_fd_sc_hd__dfxtp_1 _14409_ (.D(_02403_),
    .Q(\r1.regblock[23][6] ),
    .CLK(_01378_));
 sky130_fd_sc_hd__dfxtp_1 _14410_ (.D(_02404_),
    .Q(\r1.regblock[23][7] ),
    .CLK(_01379_));
 sky130_fd_sc_hd__dfxtp_1 _14411_ (.D(_02405_),
    .Q(\r1.regblock[23][8] ),
    .CLK(_01380_));
 sky130_fd_sc_hd__dfxtp_1 _14412_ (.D(_02406_),
    .Q(\r1.regblock[23][9] ),
    .CLK(_01381_));
 sky130_fd_sc_hd__dfxtp_1 _14413_ (.D(_02407_),
    .Q(\r1.regblock[23][10] ),
    .CLK(_01382_));
 sky130_fd_sc_hd__dfxtp_1 _14414_ (.D(_02408_),
    .Q(\r1.regblock[23][11] ),
    .CLK(_01383_));
 sky130_fd_sc_hd__dfxtp_1 _14415_ (.D(_02409_),
    .Q(\r1.regblock[23][12] ),
    .CLK(_01384_));
 sky130_fd_sc_hd__dfxtp_1 _14416_ (.D(_02410_),
    .Q(\r1.regblock[23][13] ),
    .CLK(_01385_));
 sky130_fd_sc_hd__dfxtp_1 _14417_ (.D(_02411_),
    .Q(\r1.regblock[23][14] ),
    .CLK(_01386_));
 sky130_fd_sc_hd__dfxtp_1 _14418_ (.D(_02412_),
    .Q(\r1.regblock[23][15] ),
    .CLK(_01387_));
 sky130_fd_sc_hd__dfxtp_1 _14419_ (.D(_02413_),
    .Q(\r1.regblock[23][16] ),
    .CLK(_01388_));
 sky130_fd_sc_hd__dfxtp_1 _14420_ (.D(_02414_),
    .Q(\r1.regblock[23][17] ),
    .CLK(_01389_));
 sky130_fd_sc_hd__dfxtp_1 _14421_ (.D(_02415_),
    .Q(\r1.regblock[23][18] ),
    .CLK(_01390_));
 sky130_fd_sc_hd__dfxtp_1 _14422_ (.D(_02416_),
    .Q(\r1.regblock[23][19] ),
    .CLK(_01391_));
 sky130_fd_sc_hd__dfxtp_1 _14423_ (.D(_02417_),
    .Q(\r1.regblock[23][20] ),
    .CLK(_01392_));
 sky130_fd_sc_hd__dfxtp_1 _14424_ (.D(_02418_),
    .Q(\r1.regblock[23][21] ),
    .CLK(_01393_));
 sky130_fd_sc_hd__dfxtp_1 _14425_ (.D(_02419_),
    .Q(\r1.regblock[23][22] ),
    .CLK(_01394_));
 sky130_fd_sc_hd__dfxtp_1 _14426_ (.D(_02420_),
    .Q(\r1.regblock[23][23] ),
    .CLK(_01395_));
 sky130_fd_sc_hd__dfxtp_1 _14427_ (.D(_02421_),
    .Q(\r1.regblock[23][24] ),
    .CLK(_01396_));
 sky130_fd_sc_hd__dfxtp_1 _14428_ (.D(_02422_),
    .Q(\r1.regblock[23][25] ),
    .CLK(_01397_));
 sky130_fd_sc_hd__dfxtp_1 _14429_ (.D(_02423_),
    .Q(\r1.regblock[23][26] ),
    .CLK(_01398_));
 sky130_fd_sc_hd__dfxtp_1 _14430_ (.D(_02424_),
    .Q(\r1.regblock[23][27] ),
    .CLK(_01399_));
 sky130_fd_sc_hd__dfxtp_1 _14431_ (.D(_02425_),
    .Q(\r1.regblock[23][28] ),
    .CLK(_01400_));
 sky130_fd_sc_hd__dfxtp_1 _14432_ (.D(_02426_),
    .Q(\r1.regblock[23][29] ),
    .CLK(_01401_));
 sky130_fd_sc_hd__dfxtp_1 _14433_ (.D(_02427_),
    .Q(\r1.regblock[23][30] ),
    .CLK(_01402_));
 sky130_fd_sc_hd__dfxtp_1 _14434_ (.D(_02428_),
    .Q(\r1.regblock[23][31] ),
    .CLK(_01403_));
 sky130_fd_sc_hd__dfxtp_1 _14435_ (.D(_02429_),
    .Q(\r1.regblock[22][0] ),
    .CLK(_01404_));
 sky130_fd_sc_hd__dfxtp_1 _14436_ (.D(_02430_),
    .Q(\r1.regblock[22][1] ),
    .CLK(_01405_));
 sky130_fd_sc_hd__dfxtp_1 _14437_ (.D(_02431_),
    .Q(\r1.regblock[22][2] ),
    .CLK(_01406_));
 sky130_fd_sc_hd__dfxtp_1 _14438_ (.D(_02432_),
    .Q(\r1.regblock[22][3] ),
    .CLK(_01407_));
 sky130_fd_sc_hd__dfxtp_1 _14439_ (.D(_02433_),
    .Q(\r1.regblock[22][4] ),
    .CLK(_01408_));
 sky130_fd_sc_hd__dfxtp_1 _14440_ (.D(_02434_),
    .Q(\r1.regblock[22][5] ),
    .CLK(_01409_));
 sky130_fd_sc_hd__dfxtp_1 _14441_ (.D(_02435_),
    .Q(\r1.regblock[22][6] ),
    .CLK(_01410_));
 sky130_fd_sc_hd__dfxtp_1 _14442_ (.D(_02436_),
    .Q(\r1.regblock[22][7] ),
    .CLK(_01411_));
 sky130_fd_sc_hd__dfxtp_1 _14443_ (.D(_02437_),
    .Q(\r1.regblock[22][8] ),
    .CLK(_01412_));
 sky130_fd_sc_hd__dfxtp_1 _14444_ (.D(_02438_),
    .Q(\r1.regblock[22][9] ),
    .CLK(_01413_));
 sky130_fd_sc_hd__dfxtp_1 _14445_ (.D(_02439_),
    .Q(\r1.regblock[22][10] ),
    .CLK(_01414_));
 sky130_fd_sc_hd__dfxtp_1 _14446_ (.D(_02440_),
    .Q(\r1.regblock[22][11] ),
    .CLK(_01415_));
 sky130_fd_sc_hd__dfxtp_1 _14447_ (.D(_02441_),
    .Q(\r1.regblock[22][12] ),
    .CLK(_01416_));
 sky130_fd_sc_hd__dfxtp_1 _14448_ (.D(_02442_),
    .Q(\r1.regblock[22][13] ),
    .CLK(_01417_));
 sky130_fd_sc_hd__dfxtp_1 _14449_ (.D(_02443_),
    .Q(\r1.regblock[22][14] ),
    .CLK(_01418_));
 sky130_fd_sc_hd__dfxtp_1 _14450_ (.D(_02444_),
    .Q(\r1.regblock[22][15] ),
    .CLK(_01419_));
 sky130_fd_sc_hd__dfxtp_1 _14451_ (.D(_02445_),
    .Q(\r1.regblock[22][16] ),
    .CLK(_01420_));
 sky130_fd_sc_hd__dfxtp_1 _14452_ (.D(_02446_),
    .Q(\r1.regblock[22][17] ),
    .CLK(_01421_));
 sky130_fd_sc_hd__dfxtp_1 _14453_ (.D(_02447_),
    .Q(\r1.regblock[22][18] ),
    .CLK(_01422_));
 sky130_fd_sc_hd__dfxtp_1 _14454_ (.D(_02448_),
    .Q(\r1.regblock[22][19] ),
    .CLK(_01423_));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.D(_02449_),
    .Q(\r1.regblock[22][20] ),
    .CLK(_01424_));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.D(_02450_),
    .Q(\r1.regblock[22][21] ),
    .CLK(_01425_));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.D(_02451_),
    .Q(\r1.regblock[22][22] ),
    .CLK(_01426_));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.D(_02452_),
    .Q(\r1.regblock[22][23] ),
    .CLK(_01427_));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.D(_02453_),
    .Q(\r1.regblock[22][24] ),
    .CLK(_01428_));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.D(_02454_),
    .Q(\r1.regblock[22][25] ),
    .CLK(_01429_));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.D(_02455_),
    .Q(\r1.regblock[22][26] ),
    .CLK(_01430_));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.D(_02456_),
    .Q(\r1.regblock[22][27] ),
    .CLK(_01431_));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.D(_02457_),
    .Q(\r1.regblock[22][28] ),
    .CLK(_01432_));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.D(_02458_),
    .Q(\r1.regblock[22][29] ),
    .CLK(_01433_));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.D(_02459_),
    .Q(\r1.regblock[22][30] ),
    .CLK(_01434_));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.D(_02460_),
    .Q(\r1.regblock[22][31] ),
    .CLK(_01435_));
 sky130_fd_sc_hd__dfxtp_1 _14467_ (.D(_02461_),
    .Q(\r1.regblock[21][0] ),
    .CLK(_01436_));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.D(_02462_),
    .Q(\r1.regblock[21][1] ),
    .CLK(_01437_));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.D(_02463_),
    .Q(\r1.regblock[21][2] ),
    .CLK(_01438_));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.D(_02464_),
    .Q(\r1.regblock[21][3] ),
    .CLK(_01439_));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.D(_02465_),
    .Q(\r1.regblock[21][4] ),
    .CLK(_01440_));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.D(_02466_),
    .Q(\r1.regblock[21][5] ),
    .CLK(_01441_));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.D(_02467_),
    .Q(\r1.regblock[21][6] ),
    .CLK(_01442_));
 sky130_fd_sc_hd__dfxtp_1 _14474_ (.D(_02468_),
    .Q(\r1.regblock[21][7] ),
    .CLK(_01443_));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.D(_02469_),
    .Q(\r1.regblock[21][8] ),
    .CLK(_01444_));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.D(_02470_),
    .Q(\r1.regblock[21][9] ),
    .CLK(_01445_));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.D(_02471_),
    .Q(\r1.regblock[21][10] ),
    .CLK(_01446_));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.D(_02472_),
    .Q(\r1.regblock[21][11] ),
    .CLK(_01447_));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.D(_02473_),
    .Q(\r1.regblock[21][12] ),
    .CLK(_01448_));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.D(_02474_),
    .Q(\r1.regblock[21][13] ),
    .CLK(_01449_));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.D(_02475_),
    .Q(\r1.regblock[21][14] ),
    .CLK(_01450_));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.D(_02476_),
    .Q(\r1.regblock[21][15] ),
    .CLK(_01451_));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.D(_02477_),
    .Q(\r1.regblock[21][16] ),
    .CLK(_01452_));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.D(_02478_),
    .Q(\r1.regblock[21][17] ),
    .CLK(_01453_));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.D(_02479_),
    .Q(\r1.regblock[21][18] ),
    .CLK(_01454_));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.D(_02480_),
    .Q(\r1.regblock[21][19] ),
    .CLK(_01455_));
 sky130_fd_sc_hd__dfxtp_1 _14487_ (.D(_02481_),
    .Q(\r1.regblock[21][20] ),
    .CLK(_01456_));
 sky130_fd_sc_hd__dfxtp_1 _14488_ (.D(_02482_),
    .Q(\r1.regblock[21][21] ),
    .CLK(_01457_));
 sky130_fd_sc_hd__dfxtp_1 _14489_ (.D(_02483_),
    .Q(\r1.regblock[21][22] ),
    .CLK(_01458_));
 sky130_fd_sc_hd__dfxtp_1 _14490_ (.D(_02484_),
    .Q(\r1.regblock[21][23] ),
    .CLK(_01459_));
 sky130_fd_sc_hd__dfxtp_1 _14491_ (.D(_02485_),
    .Q(\r1.regblock[21][24] ),
    .CLK(_01460_));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.D(_02486_),
    .Q(\r1.regblock[21][25] ),
    .CLK(_01461_));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.D(_02487_),
    .Q(\r1.regblock[21][26] ),
    .CLK(_01462_));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.D(_02488_),
    .Q(\r1.regblock[21][27] ),
    .CLK(_01463_));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.D(_02489_),
    .Q(\r1.regblock[21][28] ),
    .CLK(_01464_));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.D(_02490_),
    .Q(\r1.regblock[21][29] ),
    .CLK(_01465_));
 sky130_fd_sc_hd__dfxtp_1 _14497_ (.D(_02491_),
    .Q(\r1.regblock[21][30] ),
    .CLK(_01466_));
 sky130_fd_sc_hd__dfxtp_1 _14498_ (.D(_02492_),
    .Q(\r1.regblock[21][31] ),
    .CLK(_01467_));
 sky130_fd_sc_hd__dfxtp_1 _14499_ (.D(_02493_),
    .Q(\r1.regblock[20][0] ),
    .CLK(_01468_));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.D(_02494_),
    .Q(\r1.regblock[20][1] ),
    .CLK(_01469_));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.D(_02495_),
    .Q(\r1.regblock[20][2] ),
    .CLK(_01470_));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.D(_02496_),
    .Q(\r1.regblock[20][3] ),
    .CLK(_01471_));
 sky130_fd_sc_hd__dfxtp_1 _14503_ (.D(_02497_),
    .Q(\r1.regblock[20][4] ),
    .CLK(_01472_));
 sky130_fd_sc_hd__dfxtp_1 _14504_ (.D(_02498_),
    .Q(\r1.regblock[20][5] ),
    .CLK(_01473_));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.D(_02499_),
    .Q(\r1.regblock[20][6] ),
    .CLK(_01474_));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.D(_02500_),
    .Q(\r1.regblock[20][7] ),
    .CLK(_01475_));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.D(_02501_),
    .Q(\r1.regblock[20][8] ),
    .CLK(_01476_));
 sky130_fd_sc_hd__dfxtp_1 _14508_ (.D(_02502_),
    .Q(\r1.regblock[20][9] ),
    .CLK(_01477_));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.D(_02503_),
    .Q(\r1.regblock[20][10] ),
    .CLK(_01478_));
 sky130_fd_sc_hd__dfxtp_1 _14510_ (.D(_02504_),
    .Q(\r1.regblock[20][11] ),
    .CLK(_01479_));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.D(_02505_),
    .Q(\r1.regblock[20][12] ),
    .CLK(_01480_));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.D(_02506_),
    .Q(\r1.regblock[20][13] ),
    .CLK(_01481_));
 sky130_fd_sc_hd__dfxtp_1 _14513_ (.D(_02507_),
    .Q(\r1.regblock[20][14] ),
    .CLK(_01482_));
 sky130_fd_sc_hd__dfxtp_1 _14514_ (.D(_02508_),
    .Q(\r1.regblock[20][15] ),
    .CLK(_01483_));
 sky130_fd_sc_hd__dfxtp_1 _14515_ (.D(_02509_),
    .Q(\r1.regblock[20][16] ),
    .CLK(_01484_));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.D(_02510_),
    .Q(\r1.regblock[20][17] ),
    .CLK(_01485_));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.D(_02511_),
    .Q(\r1.regblock[20][18] ),
    .CLK(_01486_));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.D(_02512_),
    .Q(\r1.regblock[20][19] ),
    .CLK(_01487_));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.D(_02513_),
    .Q(\r1.regblock[20][20] ),
    .CLK(_01488_));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.D(_02514_),
    .Q(\r1.regblock[20][21] ),
    .CLK(_01489_));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.D(_02515_),
    .Q(\r1.regblock[20][22] ),
    .CLK(_01490_));
 sky130_fd_sc_hd__dfxtp_1 _14522_ (.D(_02516_),
    .Q(\r1.regblock[20][23] ),
    .CLK(_01491_));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.D(_02517_),
    .Q(\r1.regblock[20][24] ),
    .CLK(_01492_));
 sky130_fd_sc_hd__dfxtp_1 _14524_ (.D(_02518_),
    .Q(\r1.regblock[20][25] ),
    .CLK(_01493_));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.D(_02519_),
    .Q(\r1.regblock[20][26] ),
    .CLK(_01494_));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.D(_02520_),
    .Q(\r1.regblock[20][27] ),
    .CLK(_01495_));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.D(_02521_),
    .Q(\r1.regblock[20][28] ),
    .CLK(_01496_));
 sky130_fd_sc_hd__dfxtp_1 _14528_ (.D(_02522_),
    .Q(\r1.regblock[20][29] ),
    .CLK(_01497_));
 sky130_fd_sc_hd__dfxtp_1 _14529_ (.D(_02523_),
    .Q(\r1.regblock[20][30] ),
    .CLK(_01498_));
 sky130_fd_sc_hd__dfxtp_1 _14530_ (.D(_02524_),
    .Q(\r1.regblock[20][31] ),
    .CLK(_01499_));
 sky130_fd_sc_hd__dfxtp_1 _14531_ (.D(_02525_),
    .Q(\r1.regblock[1][0] ),
    .CLK(_01500_));
 sky130_fd_sc_hd__dfxtp_1 _14532_ (.D(_02526_),
    .Q(\r1.regblock[1][1] ),
    .CLK(_01501_));
 sky130_fd_sc_hd__dfxtp_1 _14533_ (.D(_02527_),
    .Q(\r1.regblock[1][2] ),
    .CLK(_01502_));
 sky130_fd_sc_hd__dfxtp_1 _14534_ (.D(_02528_),
    .Q(\r1.regblock[1][3] ),
    .CLK(_01503_));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.D(_02529_),
    .Q(\r1.regblock[1][4] ),
    .CLK(_01504_));
 sky130_fd_sc_hd__dfxtp_1 _14536_ (.D(_02530_),
    .Q(\r1.regblock[1][5] ),
    .CLK(_01505_));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.D(_02531_),
    .Q(\r1.regblock[1][6] ),
    .CLK(_01506_));
 sky130_fd_sc_hd__dfxtp_1 _14538_ (.D(_02532_),
    .Q(\r1.regblock[1][7] ),
    .CLK(_01507_));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.D(_02533_),
    .Q(\r1.regblock[1][8] ),
    .CLK(_01508_));
 sky130_fd_sc_hd__dfxtp_1 _14540_ (.D(_02534_),
    .Q(\r1.regblock[1][9] ),
    .CLK(_01509_));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.D(_02535_),
    .Q(\r1.regblock[1][10] ),
    .CLK(_01510_));
 sky130_fd_sc_hd__dfxtp_1 _14542_ (.D(_02536_),
    .Q(\r1.regblock[1][11] ),
    .CLK(_01511_));
 sky130_fd_sc_hd__dfxtp_1 _14543_ (.D(_02537_),
    .Q(\r1.regblock[1][12] ),
    .CLK(_01512_));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.D(_02538_),
    .Q(\r1.regblock[1][13] ),
    .CLK(_01513_));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.D(_02539_),
    .Q(\r1.regblock[1][14] ),
    .CLK(_01514_));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.D(_02540_),
    .Q(\r1.regblock[1][15] ),
    .CLK(_01515_));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.D(_02541_),
    .Q(\r1.regblock[1][16] ),
    .CLK(_01516_));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.D(_02542_),
    .Q(\r1.regblock[1][17] ),
    .CLK(_01517_));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.D(_02543_),
    .Q(\r1.regblock[1][18] ),
    .CLK(_01518_));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.D(_02544_),
    .Q(\r1.regblock[1][19] ),
    .CLK(_01519_));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.D(_02545_),
    .Q(\r1.regblock[1][20] ),
    .CLK(_01520_));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.D(_02546_),
    .Q(\r1.regblock[1][21] ),
    .CLK(_01521_));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.D(_02547_),
    .Q(\r1.regblock[1][22] ),
    .CLK(_01522_));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.D(_02548_),
    .Q(\r1.regblock[1][23] ),
    .CLK(_01523_));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.D(_02549_),
    .Q(\r1.regblock[1][24] ),
    .CLK(_01524_));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.D(_02550_),
    .Q(\r1.regblock[1][25] ),
    .CLK(_01525_));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.D(_02551_),
    .Q(\r1.regblock[1][26] ),
    .CLK(_01526_));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.D(_02552_),
    .Q(\r1.regblock[1][27] ),
    .CLK(_01527_));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.D(_02553_),
    .Q(\r1.regblock[1][28] ),
    .CLK(_01528_));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.D(_02554_),
    .Q(\r1.regblock[1][29] ),
    .CLK(_01529_));
 sky130_fd_sc_hd__dfxtp_1 _14561_ (.D(_02555_),
    .Q(\r1.regblock[1][30] ),
    .CLK(_01530_));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.D(_02556_),
    .Q(\r1.regblock[1][31] ),
    .CLK(_01531_));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.D(_02557_),
    .Q(\r1.regblock[18][0] ),
    .CLK(_01532_));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.D(_02558_),
    .Q(\r1.regblock[18][1] ),
    .CLK(_01533_));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.D(_02559_),
    .Q(\r1.regblock[18][2] ),
    .CLK(_01534_));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.D(_02560_),
    .Q(\r1.regblock[18][3] ),
    .CLK(_01535_));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.D(_02561_),
    .Q(\r1.regblock[18][4] ),
    .CLK(_01536_));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.D(_02562_),
    .Q(\r1.regblock[18][5] ),
    .CLK(_01537_));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.D(_02563_),
    .Q(\r1.regblock[18][6] ),
    .CLK(_01538_));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.D(_02564_),
    .Q(\r1.regblock[18][7] ),
    .CLK(_01539_));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.D(_02565_),
    .Q(\r1.regblock[18][8] ),
    .CLK(_01540_));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.D(_02566_),
    .Q(\r1.regblock[18][9] ),
    .CLK(_01541_));
 sky130_fd_sc_hd__dfxtp_1 _14573_ (.D(_02567_),
    .Q(\r1.regblock[18][10] ),
    .CLK(_01542_));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.D(_02568_),
    .Q(\r1.regblock[18][11] ),
    .CLK(_01543_));
 sky130_fd_sc_hd__dfxtp_1 _14575_ (.D(_02569_),
    .Q(\r1.regblock[18][12] ),
    .CLK(_01544_));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.D(_02570_),
    .Q(\r1.regblock[18][13] ),
    .CLK(_01545_));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.D(_02571_),
    .Q(\r1.regblock[18][14] ),
    .CLK(_01546_));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.D(_02572_),
    .Q(\r1.regblock[18][15] ),
    .CLK(_01547_));
 sky130_fd_sc_hd__dfxtp_1 _14579_ (.D(_02573_),
    .Q(\r1.regblock[18][16] ),
    .CLK(_01548_));
 sky130_fd_sc_hd__dfxtp_1 _14580_ (.D(_02574_),
    .Q(\r1.regblock[18][17] ),
    .CLK(_01549_));
 sky130_fd_sc_hd__dfxtp_1 _14581_ (.D(_02575_),
    .Q(\r1.regblock[18][18] ),
    .CLK(_01550_));
 sky130_fd_sc_hd__dfxtp_1 _14582_ (.D(_02576_),
    .Q(\r1.regblock[18][19] ),
    .CLK(_01551_));
 sky130_fd_sc_hd__dfxtp_1 _14583_ (.D(_02577_),
    .Q(\r1.regblock[18][20] ),
    .CLK(_01552_));
 sky130_fd_sc_hd__dfxtp_1 _14584_ (.D(_02578_),
    .Q(\r1.regblock[18][21] ),
    .CLK(_01553_));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.D(_02579_),
    .Q(\r1.regblock[18][22] ),
    .CLK(_01554_));
 sky130_fd_sc_hd__dfxtp_1 _14586_ (.D(_02580_),
    .Q(\r1.regblock[18][23] ),
    .CLK(_01555_));
 sky130_fd_sc_hd__dfxtp_1 _14587_ (.D(_02581_),
    .Q(\r1.regblock[18][24] ),
    .CLK(_01556_));
 sky130_fd_sc_hd__dfxtp_1 _14588_ (.D(_02582_),
    .Q(\r1.regblock[18][25] ),
    .CLK(_01557_));
 sky130_fd_sc_hd__dfxtp_1 _14589_ (.D(_02583_),
    .Q(\r1.regblock[18][26] ),
    .CLK(_01558_));
 sky130_fd_sc_hd__dfxtp_1 _14590_ (.D(_02584_),
    .Q(\r1.regblock[18][27] ),
    .CLK(_01559_));
 sky130_fd_sc_hd__dfxtp_1 _14591_ (.D(_02585_),
    .Q(\r1.regblock[18][28] ),
    .CLK(_01560_));
 sky130_fd_sc_hd__dfxtp_1 _14592_ (.D(_02586_),
    .Q(\r1.regblock[18][29] ),
    .CLK(_01561_));
 sky130_fd_sc_hd__dfxtp_1 _14593_ (.D(_02587_),
    .Q(\r1.regblock[18][30] ),
    .CLK(_01562_));
 sky130_fd_sc_hd__dfxtp_1 _14594_ (.D(_02588_),
    .Q(\r1.regblock[18][31] ),
    .CLK(_01563_));
 sky130_fd_sc_hd__dfxtp_1 _14595_ (.D(_02589_),
    .Q(\r1.regblock[17][0] ),
    .CLK(_01564_));
 sky130_fd_sc_hd__dfxtp_1 _14596_ (.D(_02590_),
    .Q(\r1.regblock[17][1] ),
    .CLK(_01565_));
 sky130_fd_sc_hd__dfxtp_1 _14597_ (.D(_02591_),
    .Q(\r1.regblock[17][2] ),
    .CLK(_01566_));
 sky130_fd_sc_hd__dfxtp_1 _14598_ (.D(_02592_),
    .Q(\r1.regblock[17][3] ),
    .CLK(_01567_));
 sky130_fd_sc_hd__dfxtp_1 _14599_ (.D(_02593_),
    .Q(\r1.regblock[17][4] ),
    .CLK(_01568_));
 sky130_fd_sc_hd__dfxtp_1 _14600_ (.D(_02594_),
    .Q(\r1.regblock[17][5] ),
    .CLK(_01569_));
 sky130_fd_sc_hd__dfxtp_1 _14601_ (.D(_02595_),
    .Q(\r1.regblock[17][6] ),
    .CLK(_01570_));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.D(_02596_),
    .Q(\r1.regblock[17][7] ),
    .CLK(_01571_));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.D(_02597_),
    .Q(\r1.regblock[17][8] ),
    .CLK(_01572_));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.D(_02598_),
    .Q(\r1.regblock[17][9] ),
    .CLK(_01573_));
 sky130_fd_sc_hd__dfxtp_1 _14605_ (.D(_02599_),
    .Q(\r1.regblock[17][10] ),
    .CLK(_01574_));
 sky130_fd_sc_hd__dfxtp_1 _14606_ (.D(_02600_),
    .Q(\r1.regblock[17][11] ),
    .CLK(_01575_));
 sky130_fd_sc_hd__dfxtp_1 _14607_ (.D(_02601_),
    .Q(\r1.regblock[17][12] ),
    .CLK(_01576_));
 sky130_fd_sc_hd__dfxtp_1 _14608_ (.D(_02602_),
    .Q(\r1.regblock[17][13] ),
    .CLK(_01577_));
 sky130_fd_sc_hd__dfxtp_1 _14609_ (.D(_02603_),
    .Q(\r1.regblock[17][14] ),
    .CLK(_01578_));
 sky130_fd_sc_hd__dfxtp_1 _14610_ (.D(_02604_),
    .Q(\r1.regblock[17][15] ),
    .CLK(_01579_));
 sky130_fd_sc_hd__dfxtp_1 _14611_ (.D(_02605_),
    .Q(\r1.regblock[17][16] ),
    .CLK(_01580_));
 sky130_fd_sc_hd__dfxtp_1 _14612_ (.D(_02606_),
    .Q(\r1.regblock[17][17] ),
    .CLK(_01581_));
 sky130_fd_sc_hd__dfxtp_1 _14613_ (.D(_02607_),
    .Q(\r1.regblock[17][18] ),
    .CLK(_01582_));
 sky130_fd_sc_hd__dfxtp_1 _14614_ (.D(_02608_),
    .Q(\r1.regblock[17][19] ),
    .CLK(_01583_));
 sky130_fd_sc_hd__dfxtp_1 _14615_ (.D(_02609_),
    .Q(\r1.regblock[17][20] ),
    .CLK(_01584_));
 sky130_fd_sc_hd__dfxtp_1 _14616_ (.D(_02610_),
    .Q(\r1.regblock[17][21] ),
    .CLK(_01585_));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.D(_02611_),
    .Q(\r1.regblock[17][22] ),
    .CLK(_01586_));
 sky130_fd_sc_hd__dfxtp_1 _14618_ (.D(_02612_),
    .Q(\r1.regblock[17][23] ),
    .CLK(_01587_));
 sky130_fd_sc_hd__dfxtp_1 _14619_ (.D(_02613_),
    .Q(\r1.regblock[17][24] ),
    .CLK(_01588_));
 sky130_fd_sc_hd__dfxtp_1 _14620_ (.D(_02614_),
    .Q(\r1.regblock[17][25] ),
    .CLK(_01589_));
 sky130_fd_sc_hd__dfxtp_1 _14621_ (.D(_02615_),
    .Q(\r1.regblock[17][26] ),
    .CLK(_01590_));
 sky130_fd_sc_hd__dfxtp_1 _14622_ (.D(_02616_),
    .Q(\r1.regblock[17][27] ),
    .CLK(_01591_));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.D(_02617_),
    .Q(\r1.regblock[17][28] ),
    .CLK(_01592_));
 sky130_fd_sc_hd__dfxtp_1 _14624_ (.D(_02618_),
    .Q(\r1.regblock[17][29] ),
    .CLK(_01593_));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.D(_02619_),
    .Q(\r1.regblock[17][30] ),
    .CLK(_01594_));
 sky130_fd_sc_hd__dfxtp_1 _14626_ (.D(_02620_),
    .Q(\r1.regblock[17][31] ),
    .CLK(_01595_));
 sky130_fd_sc_hd__dfxtp_1 _14627_ (.D(_02621_),
    .Q(\r1.regblock[16][0] ),
    .CLK(_01596_));
 sky130_fd_sc_hd__dfxtp_1 _14628_ (.D(_02622_),
    .Q(\r1.regblock[16][1] ),
    .CLK(_01597_));
 sky130_fd_sc_hd__dfxtp_1 _14629_ (.D(_02623_),
    .Q(\r1.regblock[16][2] ),
    .CLK(_01598_));
 sky130_fd_sc_hd__dfxtp_1 _14630_ (.D(_02624_),
    .Q(\r1.regblock[16][3] ),
    .CLK(_01599_));
 sky130_fd_sc_hd__dfxtp_1 _14631_ (.D(_02625_),
    .Q(\r1.regblock[16][4] ),
    .CLK(_01600_));
 sky130_fd_sc_hd__dfxtp_1 _14632_ (.D(_02626_),
    .Q(\r1.regblock[16][5] ),
    .CLK(_01601_));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.D(_02627_),
    .Q(\r1.regblock[16][6] ),
    .CLK(_01602_));
 sky130_fd_sc_hd__dfxtp_1 _14634_ (.D(_02628_),
    .Q(\r1.regblock[16][7] ),
    .CLK(_01603_));
 sky130_fd_sc_hd__dfxtp_1 _14635_ (.D(_02629_),
    .Q(\r1.regblock[16][8] ),
    .CLK(_01604_));
 sky130_fd_sc_hd__dfxtp_1 _14636_ (.D(_02630_),
    .Q(\r1.regblock[16][9] ),
    .CLK(_01605_));
 sky130_fd_sc_hd__dfxtp_1 _14637_ (.D(_02631_),
    .Q(\r1.regblock[16][10] ),
    .CLK(_01606_));
 sky130_fd_sc_hd__dfxtp_1 _14638_ (.D(_02632_),
    .Q(\r1.regblock[16][11] ),
    .CLK(_01607_));
 sky130_fd_sc_hd__dfxtp_1 _14639_ (.D(_02633_),
    .Q(\r1.regblock[16][12] ),
    .CLK(_01608_));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.D(_02634_),
    .Q(\r1.regblock[16][13] ),
    .CLK(_01609_));
 sky130_fd_sc_hd__dfxtp_1 _14641_ (.D(_02635_),
    .Q(\r1.regblock[16][14] ),
    .CLK(_01610_));
 sky130_fd_sc_hd__dfxtp_1 _14642_ (.D(_02636_),
    .Q(\r1.regblock[16][15] ),
    .CLK(_01611_));
 sky130_fd_sc_hd__dfxtp_1 _14643_ (.D(_02637_),
    .Q(\r1.regblock[16][16] ),
    .CLK(_01612_));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.D(_02638_),
    .Q(\r1.regblock[16][17] ),
    .CLK(_01613_));
 sky130_fd_sc_hd__dfxtp_1 _14645_ (.D(_02639_),
    .Q(\r1.regblock[16][18] ),
    .CLK(_01614_));
 sky130_fd_sc_hd__dfxtp_1 _14646_ (.D(_02640_),
    .Q(\r1.regblock[16][19] ),
    .CLK(_01615_));
 sky130_fd_sc_hd__dfxtp_1 _14647_ (.D(_02641_),
    .Q(\r1.regblock[16][20] ),
    .CLK(_01616_));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.D(_02642_),
    .Q(\r1.regblock[16][21] ),
    .CLK(_01617_));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.D(_02643_),
    .Q(\r1.regblock[16][22] ),
    .CLK(_01618_));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.D(_02644_),
    .Q(\r1.regblock[16][23] ),
    .CLK(_01619_));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.D(_02645_),
    .Q(\r1.regblock[16][24] ),
    .CLK(_01620_));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.D(_02646_),
    .Q(\r1.regblock[16][25] ),
    .CLK(_01621_));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.D(_02647_),
    .Q(\r1.regblock[16][26] ),
    .CLK(_01622_));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.D(_02648_),
    .Q(\r1.regblock[16][27] ),
    .CLK(_01623_));
 sky130_fd_sc_hd__dfxtp_1 _14655_ (.D(_02649_),
    .Q(\r1.regblock[16][28] ),
    .CLK(_01624_));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.D(_02650_),
    .Q(\r1.regblock[16][29] ),
    .CLK(_01625_));
 sky130_fd_sc_hd__dfxtp_1 _14657_ (.D(_02651_),
    .Q(\r1.regblock[16][30] ),
    .CLK(_01626_));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.D(_02652_),
    .Q(\r1.regblock[16][31] ),
    .CLK(_01627_));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.D(_02653_),
    .Q(\r1.regblock[4][0] ),
    .CLK(_01628_));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.D(_02654_),
    .Q(\r1.regblock[4][1] ),
    .CLK(_01629_));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.D(_02655_),
    .Q(\r1.regblock[4][2] ),
    .CLK(_01630_));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.D(_02656_),
    .Q(\r1.regblock[4][3] ),
    .CLK(_01631_));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.D(_02657_),
    .Q(\r1.regblock[4][4] ),
    .CLK(_01632_));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.D(_02658_),
    .Q(\r1.regblock[4][5] ),
    .CLK(_01633_));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.D(_02659_),
    .Q(\r1.regblock[4][6] ),
    .CLK(_01634_));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.D(_02660_),
    .Q(\r1.regblock[4][7] ),
    .CLK(_01635_));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.D(_02661_),
    .Q(\r1.regblock[4][8] ),
    .CLK(_01636_));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.D(_02662_),
    .Q(\r1.regblock[4][9] ),
    .CLK(_01637_));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.D(_02663_),
    .Q(\r1.regblock[4][10] ),
    .CLK(_01638_));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.D(_02664_),
    .Q(\r1.regblock[4][11] ),
    .CLK(_01639_));
 sky130_fd_sc_hd__dfxtp_1 _14671_ (.D(_02665_),
    .Q(\r1.regblock[4][12] ),
    .CLK(_01640_));
 sky130_fd_sc_hd__dfxtp_1 _14672_ (.D(_02666_),
    .Q(\r1.regblock[4][13] ),
    .CLK(_01641_));
 sky130_fd_sc_hd__dfxtp_1 _14673_ (.D(_02667_),
    .Q(\r1.regblock[4][14] ),
    .CLK(_01642_));
 sky130_fd_sc_hd__dfxtp_1 _14674_ (.D(_02668_),
    .Q(\r1.regblock[4][15] ),
    .CLK(_01643_));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.D(_02669_),
    .Q(\r1.regblock[4][16] ),
    .CLK(_01644_));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.D(_02670_),
    .Q(\r1.regblock[4][17] ),
    .CLK(_01645_));
 sky130_fd_sc_hd__dfxtp_1 _14677_ (.D(_02671_),
    .Q(\r1.regblock[4][18] ),
    .CLK(_01646_));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.D(_02672_),
    .Q(\r1.regblock[4][19] ),
    .CLK(_01647_));
 sky130_fd_sc_hd__dfxtp_1 _14679_ (.D(_02673_),
    .Q(\r1.regblock[4][20] ),
    .CLK(_01648_));
 sky130_fd_sc_hd__dfxtp_1 _14680_ (.D(_02674_),
    .Q(\r1.regblock[4][21] ),
    .CLK(_01649_));
 sky130_fd_sc_hd__dfxtp_1 _14681_ (.D(_02675_),
    .Q(\r1.regblock[4][22] ),
    .CLK(_01650_));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.D(_02676_),
    .Q(\r1.regblock[4][23] ),
    .CLK(_01651_));
 sky130_fd_sc_hd__dfxtp_1 _14683_ (.D(_02677_),
    .Q(\r1.regblock[4][24] ),
    .CLK(_01652_));
 sky130_fd_sc_hd__dfxtp_1 _14684_ (.D(_02678_),
    .Q(\r1.regblock[4][25] ),
    .CLK(_01653_));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.D(_02679_),
    .Q(\r1.regblock[4][26] ),
    .CLK(_01654_));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.D(_02680_),
    .Q(\r1.regblock[4][27] ),
    .CLK(_01655_));
 sky130_fd_sc_hd__dfxtp_1 _14687_ (.D(_02681_),
    .Q(\r1.regblock[4][28] ),
    .CLK(_01656_));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.D(_02682_),
    .Q(\r1.regblock[4][29] ),
    .CLK(_01657_));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.D(_02683_),
    .Q(\r1.regblock[4][30] ),
    .CLK(_01658_));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.D(_02684_),
    .Q(\r1.regblock[4][31] ),
    .CLK(_01659_));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.D(_02685_),
    .Q(\r1.regblock[7][0] ),
    .CLK(_01660_));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.D(_02686_),
    .Q(\r1.regblock[7][1] ),
    .CLK(_01661_));
 sky130_fd_sc_hd__dfxtp_1 _14693_ (.D(_02687_),
    .Q(\r1.regblock[7][2] ),
    .CLK(_01662_));
 sky130_fd_sc_hd__dfxtp_1 _14694_ (.D(_02688_),
    .Q(\r1.regblock[7][3] ),
    .CLK(_01663_));
 sky130_fd_sc_hd__dfxtp_1 _14695_ (.D(_02689_),
    .Q(\r1.regblock[7][4] ),
    .CLK(_01664_));
 sky130_fd_sc_hd__dfxtp_1 _14696_ (.D(_02690_),
    .Q(\r1.regblock[7][5] ),
    .CLK(_01665_));
 sky130_fd_sc_hd__dfxtp_1 _14697_ (.D(_02691_),
    .Q(\r1.regblock[7][6] ),
    .CLK(_01666_));
 sky130_fd_sc_hd__dfxtp_1 _14698_ (.D(_02692_),
    .Q(\r1.regblock[7][7] ),
    .CLK(_01667_));
 sky130_fd_sc_hd__dfxtp_1 _14699_ (.D(_02693_),
    .Q(\r1.regblock[7][8] ),
    .CLK(_01668_));
 sky130_fd_sc_hd__dfxtp_1 _14700_ (.D(_02694_),
    .Q(\r1.regblock[7][9] ),
    .CLK(_01669_));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.D(_02695_),
    .Q(\r1.regblock[7][10] ),
    .CLK(_01670_));
 sky130_fd_sc_hd__dfxtp_1 _14702_ (.D(_02696_),
    .Q(\r1.regblock[7][11] ),
    .CLK(_01671_));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.D(_02697_),
    .Q(\r1.regblock[7][12] ),
    .CLK(_01672_));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.D(_02698_),
    .Q(\r1.regblock[7][13] ),
    .CLK(_01673_));
 sky130_fd_sc_hd__dfxtp_1 _14705_ (.D(_02699_),
    .Q(\r1.regblock[7][14] ),
    .CLK(_01674_));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.D(_02700_),
    .Q(\r1.regblock[7][15] ),
    .CLK(_01675_));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.D(_02701_),
    .Q(\r1.regblock[7][16] ),
    .CLK(_01676_));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.D(_02702_),
    .Q(\r1.regblock[7][17] ),
    .CLK(_01677_));
 sky130_fd_sc_hd__dfxtp_1 _14709_ (.D(_02703_),
    .Q(\r1.regblock[7][18] ),
    .CLK(_01678_));
 sky130_fd_sc_hd__dfxtp_1 _14710_ (.D(_02704_),
    .Q(\r1.regblock[7][19] ),
    .CLK(_01679_));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.D(_02705_),
    .Q(\r1.regblock[7][20] ),
    .CLK(_01680_));
 sky130_fd_sc_hd__dfxtp_1 _14712_ (.D(_02706_),
    .Q(\r1.regblock[7][21] ),
    .CLK(_01681_));
 sky130_fd_sc_hd__dfxtp_1 _14713_ (.D(_02707_),
    .Q(\r1.regblock[7][22] ),
    .CLK(_01682_));
 sky130_fd_sc_hd__dfxtp_1 _14714_ (.D(_02708_),
    .Q(\r1.regblock[7][23] ),
    .CLK(_01683_));
 sky130_fd_sc_hd__dfxtp_1 _14715_ (.D(_02709_),
    .Q(\r1.regblock[7][24] ),
    .CLK(_01684_));
 sky130_fd_sc_hd__dfxtp_1 _14716_ (.D(_02710_),
    .Q(\r1.regblock[7][25] ),
    .CLK(_01685_));
 sky130_fd_sc_hd__dfxtp_1 _14717_ (.D(_02711_),
    .Q(\r1.regblock[7][26] ),
    .CLK(_01686_));
 sky130_fd_sc_hd__dfxtp_1 _14718_ (.D(_02712_),
    .Q(\r1.regblock[7][27] ),
    .CLK(_01687_));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.D(_02713_),
    .Q(\r1.regblock[7][28] ),
    .CLK(_01688_));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.D(_02714_),
    .Q(\r1.regblock[7][29] ),
    .CLK(_01689_));
 sky130_fd_sc_hd__dfxtp_1 _14721_ (.D(_02715_),
    .Q(\r1.regblock[7][30] ),
    .CLK(_01690_));
 sky130_fd_sc_hd__dfxtp_1 _14722_ (.D(_02716_),
    .Q(\r1.regblock[7][31] ),
    .CLK(_01691_));
 sky130_fd_sc_hd__dfxtp_1 _14723_ (.D(_02717_),
    .Q(\r1.regblock[6][0] ),
    .CLK(_01692_));
 sky130_fd_sc_hd__dfxtp_1 _14724_ (.D(_02718_),
    .Q(\r1.regblock[6][1] ),
    .CLK(_01693_));
 sky130_fd_sc_hd__dfxtp_1 _14725_ (.D(_02719_),
    .Q(\r1.regblock[6][2] ),
    .CLK(_01694_));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.D(_02720_),
    .Q(\r1.regblock[6][3] ),
    .CLK(_01695_));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.D(_02721_),
    .Q(\r1.regblock[6][4] ),
    .CLK(_01696_));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.D(_02722_),
    .Q(\r1.regblock[6][5] ),
    .CLK(_01697_));
 sky130_fd_sc_hd__dfxtp_1 _14729_ (.D(_02723_),
    .Q(\r1.regblock[6][6] ),
    .CLK(_01698_));
 sky130_fd_sc_hd__dfxtp_1 _14730_ (.D(_02724_),
    .Q(\r1.regblock[6][7] ),
    .CLK(_01699_));
 sky130_fd_sc_hd__dfxtp_1 _14731_ (.D(_02725_),
    .Q(\r1.regblock[6][8] ),
    .CLK(_01700_));
 sky130_fd_sc_hd__dfxtp_1 _14732_ (.D(_02726_),
    .Q(\r1.regblock[6][9] ),
    .CLK(_01701_));
 sky130_fd_sc_hd__dfxtp_1 _14733_ (.D(_02727_),
    .Q(\r1.regblock[6][10] ),
    .CLK(_01702_));
 sky130_fd_sc_hd__dfxtp_1 _14734_ (.D(_02728_),
    .Q(\r1.regblock[6][11] ),
    .CLK(_01703_));
 sky130_fd_sc_hd__dfxtp_1 _14735_ (.D(_02729_),
    .Q(\r1.regblock[6][12] ),
    .CLK(_01704_));
 sky130_fd_sc_hd__dfxtp_1 _14736_ (.D(_02730_),
    .Q(\r1.regblock[6][13] ),
    .CLK(_01705_));
 sky130_fd_sc_hd__dfxtp_1 _14737_ (.D(_02731_),
    .Q(\r1.regblock[6][14] ),
    .CLK(_01706_));
 sky130_fd_sc_hd__dfxtp_1 _14738_ (.D(_02732_),
    .Q(\r1.regblock[6][15] ),
    .CLK(_01707_));
 sky130_fd_sc_hd__dfxtp_1 _14739_ (.D(_02733_),
    .Q(\r1.regblock[6][16] ),
    .CLK(_01708_));
 sky130_fd_sc_hd__dfxtp_1 _14740_ (.D(_02734_),
    .Q(\r1.regblock[6][17] ),
    .CLK(_01709_));
 sky130_fd_sc_hd__dfxtp_1 _14741_ (.D(_02735_),
    .Q(\r1.regblock[6][18] ),
    .CLK(_01710_));
 sky130_fd_sc_hd__dfxtp_1 _14742_ (.D(_02736_),
    .Q(\r1.regblock[6][19] ),
    .CLK(_01711_));
 sky130_fd_sc_hd__dfxtp_1 _14743_ (.D(_02737_),
    .Q(\r1.regblock[6][20] ),
    .CLK(_01712_));
 sky130_fd_sc_hd__dfxtp_1 _14744_ (.D(_02738_),
    .Q(\r1.regblock[6][21] ),
    .CLK(_01713_));
 sky130_fd_sc_hd__dfxtp_1 _14745_ (.D(_02739_),
    .Q(\r1.regblock[6][22] ),
    .CLK(_01714_));
 sky130_fd_sc_hd__dfxtp_1 _14746_ (.D(_02740_),
    .Q(\r1.regblock[6][23] ),
    .CLK(_01715_));
 sky130_fd_sc_hd__dfxtp_1 _14747_ (.D(_02741_),
    .Q(\r1.regblock[6][24] ),
    .CLK(_01716_));
 sky130_fd_sc_hd__dfxtp_1 _14748_ (.D(_02742_),
    .Q(\r1.regblock[6][25] ),
    .CLK(_01717_));
 sky130_fd_sc_hd__dfxtp_1 _14749_ (.D(_02743_),
    .Q(\r1.regblock[6][26] ),
    .CLK(_01718_));
 sky130_fd_sc_hd__dfxtp_1 _14750_ (.D(_02744_),
    .Q(\r1.regblock[6][27] ),
    .CLK(_01719_));
 sky130_fd_sc_hd__dfxtp_1 _14751_ (.D(_02745_),
    .Q(\r1.regblock[6][28] ),
    .CLK(_01720_));
 sky130_fd_sc_hd__dfxtp_1 _14752_ (.D(_02746_),
    .Q(\r1.regblock[6][29] ),
    .CLK(_01721_));
 sky130_fd_sc_hd__dfxtp_1 _14753_ (.D(_02747_),
    .Q(\r1.regblock[6][30] ),
    .CLK(_01722_));
 sky130_fd_sc_hd__dfxtp_1 _14754_ (.D(_02748_),
    .Q(\r1.regblock[6][31] ),
    .CLK(_01723_));
 sky130_fd_sc_hd__dfxtp_1 _14755_ (.D(_02749_),
    .Q(\r1.regblock[10][0] ),
    .CLK(_01724_));
 sky130_fd_sc_hd__dfxtp_1 _14756_ (.D(_02750_),
    .Q(\r1.regblock[10][1] ),
    .CLK(_01725_));
 sky130_fd_sc_hd__dfxtp_1 _14757_ (.D(_02751_),
    .Q(\r1.regblock[10][2] ),
    .CLK(_01726_));
 sky130_fd_sc_hd__dfxtp_1 _14758_ (.D(_02752_),
    .Q(\r1.regblock[10][3] ),
    .CLK(_01727_));
 sky130_fd_sc_hd__dfxtp_1 _14759_ (.D(_02753_),
    .Q(\r1.regblock[10][4] ),
    .CLK(_01728_));
 sky130_fd_sc_hd__dfxtp_1 _14760_ (.D(_02754_),
    .Q(\r1.regblock[10][5] ),
    .CLK(_01729_));
 sky130_fd_sc_hd__dfxtp_1 _14761_ (.D(_02755_),
    .Q(\r1.regblock[10][6] ),
    .CLK(_01730_));
 sky130_fd_sc_hd__dfxtp_1 _14762_ (.D(_02756_),
    .Q(\r1.regblock[10][7] ),
    .CLK(_01731_));
 sky130_fd_sc_hd__dfxtp_1 _14763_ (.D(_02757_),
    .Q(\r1.regblock[10][8] ),
    .CLK(_01732_));
 sky130_fd_sc_hd__dfxtp_1 _14764_ (.D(_02758_),
    .Q(\r1.regblock[10][9] ),
    .CLK(_01733_));
 sky130_fd_sc_hd__dfxtp_1 _14765_ (.D(_02759_),
    .Q(\r1.regblock[10][10] ),
    .CLK(_01734_));
 sky130_fd_sc_hd__dfxtp_1 _14766_ (.D(_02760_),
    .Q(\r1.regblock[10][11] ),
    .CLK(_01735_));
 sky130_fd_sc_hd__dfxtp_1 _14767_ (.D(_02761_),
    .Q(\r1.regblock[10][12] ),
    .CLK(_01736_));
 sky130_fd_sc_hd__dfxtp_1 _14768_ (.D(_02762_),
    .Q(\r1.regblock[10][13] ),
    .CLK(_01737_));
 sky130_fd_sc_hd__dfxtp_1 _14769_ (.D(_02763_),
    .Q(\r1.regblock[10][14] ),
    .CLK(_01738_));
 sky130_fd_sc_hd__dfxtp_1 _14770_ (.D(_02764_),
    .Q(\r1.regblock[10][15] ),
    .CLK(_01739_));
 sky130_fd_sc_hd__dfxtp_1 _14771_ (.D(_02765_),
    .Q(\r1.regblock[10][16] ),
    .CLK(_01740_));
 sky130_fd_sc_hd__dfxtp_1 _14772_ (.D(_02766_),
    .Q(\r1.regblock[10][17] ),
    .CLK(_01741_));
 sky130_fd_sc_hd__dfxtp_1 _14773_ (.D(_02767_),
    .Q(\r1.regblock[10][18] ),
    .CLK(_01742_));
 sky130_fd_sc_hd__dfxtp_1 _14774_ (.D(_02768_),
    .Q(\r1.regblock[10][19] ),
    .CLK(_01743_));
 sky130_fd_sc_hd__dfxtp_1 _14775_ (.D(_02769_),
    .Q(\r1.regblock[10][20] ),
    .CLK(_01744_));
 sky130_fd_sc_hd__dfxtp_1 _14776_ (.D(_02770_),
    .Q(\r1.regblock[10][21] ),
    .CLK(_01745_));
 sky130_fd_sc_hd__dfxtp_1 _14777_ (.D(_02771_),
    .Q(\r1.regblock[10][22] ),
    .CLK(_01746_));
 sky130_fd_sc_hd__dfxtp_1 _14778_ (.D(_02772_),
    .Q(\r1.regblock[10][23] ),
    .CLK(_01747_));
 sky130_fd_sc_hd__dfxtp_1 _14779_ (.D(_02773_),
    .Q(\r1.regblock[10][24] ),
    .CLK(_01748_));
 sky130_fd_sc_hd__dfxtp_1 _14780_ (.D(_02774_),
    .Q(\r1.regblock[10][25] ),
    .CLK(_01749_));
 sky130_fd_sc_hd__dfxtp_1 _14781_ (.D(_02775_),
    .Q(\r1.regblock[10][26] ),
    .CLK(_01750_));
 sky130_fd_sc_hd__dfxtp_1 _14782_ (.D(_02776_),
    .Q(\r1.regblock[10][27] ),
    .CLK(_01751_));
 sky130_fd_sc_hd__dfxtp_1 _14783_ (.D(_02777_),
    .Q(\r1.regblock[10][28] ),
    .CLK(_01752_));
 sky130_fd_sc_hd__dfxtp_1 _14784_ (.D(_02778_),
    .Q(\r1.regblock[10][29] ),
    .CLK(_01753_));
 sky130_fd_sc_hd__dfxtp_1 _14785_ (.D(_02779_),
    .Q(\r1.regblock[10][30] ),
    .CLK(_01754_));
 sky130_fd_sc_hd__dfxtp_1 _14786_ (.D(_02780_),
    .Q(\r1.regblock[10][31] ),
    .CLK(_01755_));
 sky130_fd_sc_hd__dfxtp_1 _14787_ (.D(_02781_),
    .Q(\r1.regblock[11][0] ),
    .CLK(_01756_));
 sky130_fd_sc_hd__dfxtp_1 _14788_ (.D(_02782_),
    .Q(\r1.regblock[11][1] ),
    .CLK(_01757_));
 sky130_fd_sc_hd__dfxtp_1 _14789_ (.D(_02783_),
    .Q(\r1.regblock[11][2] ),
    .CLK(_01758_));
 sky130_fd_sc_hd__dfxtp_1 _14790_ (.D(_02784_),
    .Q(\r1.regblock[11][3] ),
    .CLK(_01759_));
 sky130_fd_sc_hd__dfxtp_1 _14791_ (.D(_02785_),
    .Q(\r1.regblock[11][4] ),
    .CLK(_01760_));
 sky130_fd_sc_hd__dfxtp_1 _14792_ (.D(_02786_),
    .Q(\r1.regblock[11][5] ),
    .CLK(_01761_));
 sky130_fd_sc_hd__dfxtp_1 _14793_ (.D(_02787_),
    .Q(\r1.regblock[11][6] ),
    .CLK(_01762_));
 sky130_fd_sc_hd__dfxtp_1 _14794_ (.D(_02788_),
    .Q(\r1.regblock[11][7] ),
    .CLK(_01763_));
 sky130_fd_sc_hd__dfxtp_1 _14795_ (.D(_02789_),
    .Q(\r1.regblock[11][8] ),
    .CLK(_01764_));
 sky130_fd_sc_hd__dfxtp_1 _14796_ (.D(_02790_),
    .Q(\r1.regblock[11][9] ),
    .CLK(_01765_));
 sky130_fd_sc_hd__dfxtp_1 _14797_ (.D(_02791_),
    .Q(\r1.regblock[11][10] ),
    .CLK(_01766_));
 sky130_fd_sc_hd__dfxtp_1 _14798_ (.D(_02792_),
    .Q(\r1.regblock[11][11] ),
    .CLK(_01767_));
 sky130_fd_sc_hd__dfxtp_1 _14799_ (.D(_02793_),
    .Q(\r1.regblock[11][12] ),
    .CLK(_01768_));
 sky130_fd_sc_hd__dfxtp_1 _14800_ (.D(_02794_),
    .Q(\r1.regblock[11][13] ),
    .CLK(_01769_));
 sky130_fd_sc_hd__dfxtp_1 _14801_ (.D(_02795_),
    .Q(\r1.regblock[11][14] ),
    .CLK(_01770_));
 sky130_fd_sc_hd__dfxtp_1 _14802_ (.D(_02796_),
    .Q(\r1.regblock[11][15] ),
    .CLK(_01771_));
 sky130_fd_sc_hd__dfxtp_1 _14803_ (.D(_02797_),
    .Q(\r1.regblock[11][16] ),
    .CLK(_01772_));
 sky130_fd_sc_hd__dfxtp_1 _14804_ (.D(_02798_),
    .Q(\r1.regblock[11][17] ),
    .CLK(_01773_));
 sky130_fd_sc_hd__dfxtp_1 _14805_ (.D(_02799_),
    .Q(\r1.regblock[11][18] ),
    .CLK(_01774_));
 sky130_fd_sc_hd__dfxtp_1 _14806_ (.D(_02800_),
    .Q(\r1.regblock[11][19] ),
    .CLK(_01775_));
 sky130_fd_sc_hd__dfxtp_1 _14807_ (.D(_02801_),
    .Q(\r1.regblock[11][20] ),
    .CLK(_01776_));
 sky130_fd_sc_hd__dfxtp_1 _14808_ (.D(_02802_),
    .Q(\r1.regblock[11][21] ),
    .CLK(_01777_));
 sky130_fd_sc_hd__dfxtp_1 _14809_ (.D(_02803_),
    .Q(\r1.regblock[11][22] ),
    .CLK(_01778_));
 sky130_fd_sc_hd__dfxtp_1 _14810_ (.D(_02804_),
    .Q(\r1.regblock[11][23] ),
    .CLK(_01779_));
 sky130_fd_sc_hd__dfxtp_1 _14811_ (.D(_02805_),
    .Q(\r1.regblock[11][24] ),
    .CLK(_01780_));
 sky130_fd_sc_hd__dfxtp_1 _14812_ (.D(_02806_),
    .Q(\r1.regblock[11][25] ),
    .CLK(_01781_));
 sky130_fd_sc_hd__dfxtp_1 _14813_ (.D(_02807_),
    .Q(\r1.regblock[11][26] ),
    .CLK(_01782_));
 sky130_fd_sc_hd__dfxtp_1 _14814_ (.D(_02808_),
    .Q(\r1.regblock[11][27] ),
    .CLK(_01783_));
 sky130_fd_sc_hd__dfxtp_1 _14815_ (.D(_02809_),
    .Q(\r1.regblock[11][28] ),
    .CLK(_01784_));
 sky130_fd_sc_hd__dfxtp_1 _14816_ (.D(_02810_),
    .Q(\r1.regblock[11][29] ),
    .CLK(_01785_));
 sky130_fd_sc_hd__dfxtp_1 _14817_ (.D(_02811_),
    .Q(\r1.regblock[11][30] ),
    .CLK(_01786_));
 sky130_fd_sc_hd__dfxtp_1 _14818_ (.D(_02812_),
    .Q(\r1.regblock[11][31] ),
    .CLK(_01787_));
 sky130_fd_sc_hd__dfxtp_1 _14819_ (.D(_02813_),
    .Q(\r1.regblock[24][0] ),
    .CLK(_01788_));
 sky130_fd_sc_hd__dfxtp_1 _14820_ (.D(_02814_),
    .Q(\r1.regblock[24][1] ),
    .CLK(_01789_));
 sky130_fd_sc_hd__dfxtp_1 _14821_ (.D(_02815_),
    .Q(\r1.regblock[24][2] ),
    .CLK(_01790_));
 sky130_fd_sc_hd__dfxtp_1 _14822_ (.D(_02816_),
    .Q(\r1.regblock[24][3] ),
    .CLK(_01791_));
 sky130_fd_sc_hd__dfxtp_1 _14823_ (.D(_02817_),
    .Q(\r1.regblock[24][4] ),
    .CLK(_01792_));
 sky130_fd_sc_hd__dfxtp_1 _14824_ (.D(_02818_),
    .Q(\r1.regblock[24][5] ),
    .CLK(_01793_));
 sky130_fd_sc_hd__dfxtp_1 _14825_ (.D(_02819_),
    .Q(\r1.regblock[24][6] ),
    .CLK(_01794_));
 sky130_fd_sc_hd__dfxtp_1 _14826_ (.D(_02820_),
    .Q(\r1.regblock[24][7] ),
    .CLK(_01795_));
 sky130_fd_sc_hd__dfxtp_1 _14827_ (.D(_02821_),
    .Q(\r1.regblock[24][8] ),
    .CLK(_01796_));
 sky130_fd_sc_hd__dfxtp_1 _14828_ (.D(_02822_),
    .Q(\r1.regblock[24][9] ),
    .CLK(_01797_));
 sky130_fd_sc_hd__dfxtp_1 _14829_ (.D(_02823_),
    .Q(\r1.regblock[24][10] ),
    .CLK(_01798_));
 sky130_fd_sc_hd__dfxtp_1 _14830_ (.D(_02824_),
    .Q(\r1.regblock[24][11] ),
    .CLK(_01799_));
 sky130_fd_sc_hd__dfxtp_1 _14831_ (.D(_02825_),
    .Q(\r1.regblock[24][12] ),
    .CLK(_01800_));
 sky130_fd_sc_hd__dfxtp_1 _14832_ (.D(_02826_),
    .Q(\r1.regblock[24][13] ),
    .CLK(_01801_));
 sky130_fd_sc_hd__dfxtp_1 _14833_ (.D(_02827_),
    .Q(\r1.regblock[24][14] ),
    .CLK(_01802_));
 sky130_fd_sc_hd__dfxtp_1 _14834_ (.D(_02828_),
    .Q(\r1.regblock[24][15] ),
    .CLK(_01803_));
 sky130_fd_sc_hd__dfxtp_1 _14835_ (.D(_02829_),
    .Q(\r1.regblock[24][16] ),
    .CLK(_01804_));
 sky130_fd_sc_hd__dfxtp_1 _14836_ (.D(_02830_),
    .Q(\r1.regblock[24][17] ),
    .CLK(_01805_));
 sky130_fd_sc_hd__dfxtp_1 _14837_ (.D(_02831_),
    .Q(\r1.regblock[24][18] ),
    .CLK(_01806_));
 sky130_fd_sc_hd__dfxtp_1 _14838_ (.D(_02832_),
    .Q(\r1.regblock[24][19] ),
    .CLK(_01807_));
 sky130_fd_sc_hd__dfxtp_1 _14839_ (.D(_02833_),
    .Q(\r1.regblock[24][20] ),
    .CLK(_01808_));
 sky130_fd_sc_hd__dfxtp_1 _14840_ (.D(_02834_),
    .Q(\r1.regblock[24][21] ),
    .CLK(_01809_));
 sky130_fd_sc_hd__dfxtp_1 _14841_ (.D(_02835_),
    .Q(\r1.regblock[24][22] ),
    .CLK(_01810_));
 sky130_fd_sc_hd__dfxtp_1 _14842_ (.D(_02836_),
    .Q(\r1.regblock[24][23] ),
    .CLK(_01811_));
 sky130_fd_sc_hd__dfxtp_1 _14843_ (.D(_02837_),
    .Q(\r1.regblock[24][24] ),
    .CLK(_01812_));
 sky130_fd_sc_hd__dfxtp_1 _14844_ (.D(_02838_),
    .Q(\r1.regblock[24][25] ),
    .CLK(_01813_));
 sky130_fd_sc_hd__dfxtp_1 _14845_ (.D(_02839_),
    .Q(\r1.regblock[24][26] ),
    .CLK(_01814_));
 sky130_fd_sc_hd__dfxtp_1 _14846_ (.D(_02840_),
    .Q(\r1.regblock[24][27] ),
    .CLK(_01815_));
 sky130_fd_sc_hd__dfxtp_1 _14847_ (.D(_02841_),
    .Q(\r1.regblock[24][28] ),
    .CLK(_01816_));
 sky130_fd_sc_hd__dfxtp_1 _14848_ (.D(_02842_),
    .Q(\r1.regblock[24][29] ),
    .CLK(_01817_));
 sky130_fd_sc_hd__dfxtp_1 _14849_ (.D(_02843_),
    .Q(\r1.regblock[24][30] ),
    .CLK(_01818_));
 sky130_fd_sc_hd__dfxtp_1 _14850_ (.D(_02844_),
    .Q(\r1.regblock[24][31] ),
    .CLK(_01819_));
 sky130_fd_sc_hd__dfxtp_1 _14851_ (.D(_02845_),
    .Q(\r1.regblock[25][0] ),
    .CLK(_01820_));
 sky130_fd_sc_hd__dfxtp_1 _14852_ (.D(_02846_),
    .Q(\r1.regblock[25][1] ),
    .CLK(_01821_));
 sky130_fd_sc_hd__dfxtp_1 _14853_ (.D(_02847_),
    .Q(\r1.regblock[25][2] ),
    .CLK(_01822_));
 sky130_fd_sc_hd__dfxtp_1 _14854_ (.D(_02848_),
    .Q(\r1.regblock[25][3] ),
    .CLK(_01823_));
 sky130_fd_sc_hd__dfxtp_1 _14855_ (.D(_02849_),
    .Q(\r1.regblock[25][4] ),
    .CLK(_01824_));
 sky130_fd_sc_hd__dfxtp_1 _14856_ (.D(_02850_),
    .Q(\r1.regblock[25][5] ),
    .CLK(_01825_));
 sky130_fd_sc_hd__dfxtp_1 _14857_ (.D(_02851_),
    .Q(\r1.regblock[25][6] ),
    .CLK(_01826_));
 sky130_fd_sc_hd__dfxtp_1 _14858_ (.D(_02852_),
    .Q(\r1.regblock[25][7] ),
    .CLK(_01827_));
 sky130_fd_sc_hd__dfxtp_1 _14859_ (.D(_02853_),
    .Q(\r1.regblock[25][8] ),
    .CLK(_01828_));
 sky130_fd_sc_hd__dfxtp_1 _14860_ (.D(_02854_),
    .Q(\r1.regblock[25][9] ),
    .CLK(_01829_));
 sky130_fd_sc_hd__dfxtp_1 _14861_ (.D(_02855_),
    .Q(\r1.regblock[25][10] ),
    .CLK(_01830_));
 sky130_fd_sc_hd__dfxtp_1 _14862_ (.D(_02856_),
    .Q(\r1.regblock[25][11] ),
    .CLK(_01831_));
 sky130_fd_sc_hd__dfxtp_1 _14863_ (.D(_02857_),
    .Q(\r1.regblock[25][12] ),
    .CLK(_01832_));
 sky130_fd_sc_hd__dfxtp_1 _14864_ (.D(_02858_),
    .Q(\r1.regblock[25][13] ),
    .CLK(_01833_));
 sky130_fd_sc_hd__dfxtp_1 _14865_ (.D(_02859_),
    .Q(\r1.regblock[25][14] ),
    .CLK(_01834_));
 sky130_fd_sc_hd__dfxtp_1 _14866_ (.D(_02860_),
    .Q(\r1.regblock[25][15] ),
    .CLK(_01835_));
 sky130_fd_sc_hd__dfxtp_1 _14867_ (.D(_02861_),
    .Q(\r1.regblock[25][16] ),
    .CLK(_01836_));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.D(_02862_),
    .Q(\r1.regblock[25][17] ),
    .CLK(_01837_));
 sky130_fd_sc_hd__dfxtp_1 _14869_ (.D(_02863_),
    .Q(\r1.regblock[25][18] ),
    .CLK(_01838_));
 sky130_fd_sc_hd__dfxtp_1 _14870_ (.D(_02864_),
    .Q(\r1.regblock[25][19] ),
    .CLK(_01839_));
 sky130_fd_sc_hd__dfxtp_1 _14871_ (.D(_02865_),
    .Q(\r1.regblock[25][20] ),
    .CLK(_01840_));
 sky130_fd_sc_hd__dfxtp_1 _14872_ (.D(_02866_),
    .Q(\r1.regblock[25][21] ),
    .CLK(_01841_));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.D(_02867_),
    .Q(\r1.regblock[25][22] ),
    .CLK(_01842_));
 sky130_fd_sc_hd__dfxtp_1 _14874_ (.D(_02868_),
    .Q(\r1.regblock[25][23] ),
    .CLK(_01843_));
 sky130_fd_sc_hd__dfxtp_1 _14875_ (.D(_02869_),
    .Q(\r1.regblock[25][24] ),
    .CLK(_01844_));
 sky130_fd_sc_hd__dfxtp_1 _14876_ (.D(_02870_),
    .Q(\r1.regblock[25][25] ),
    .CLK(_01845_));
 sky130_fd_sc_hd__dfxtp_1 _14877_ (.D(_02871_),
    .Q(\r1.regblock[25][26] ),
    .CLK(_01846_));
 sky130_fd_sc_hd__dfxtp_1 _14878_ (.D(_02872_),
    .Q(\r1.regblock[25][27] ),
    .CLK(_01847_));
 sky130_fd_sc_hd__dfxtp_1 _14879_ (.D(_02873_),
    .Q(\r1.regblock[25][28] ),
    .CLK(_01848_));
 sky130_fd_sc_hd__dfxtp_1 _14880_ (.D(_02874_),
    .Q(\r1.regblock[25][29] ),
    .CLK(_01849_));
 sky130_fd_sc_hd__dfxtp_1 _14881_ (.D(_02875_),
    .Q(\r1.regblock[25][30] ),
    .CLK(_01850_));
 sky130_fd_sc_hd__dfxtp_1 _14882_ (.D(_02876_),
    .Q(\r1.regblock[25][31] ),
    .CLK(_01851_));
 sky130_fd_sc_hd__dfxtp_1 _14883_ (.D(_02877_),
    .Q(\r1.regblock[26][0] ),
    .CLK(_01852_));
 sky130_fd_sc_hd__dfxtp_1 _14884_ (.D(_02878_),
    .Q(\r1.regblock[26][1] ),
    .CLK(_01853_));
 sky130_fd_sc_hd__dfxtp_1 _14885_ (.D(_02879_),
    .Q(\r1.regblock[26][2] ),
    .CLK(_01854_));
 sky130_fd_sc_hd__dfxtp_1 _14886_ (.D(_02880_),
    .Q(\r1.regblock[26][3] ),
    .CLK(_01855_));
 sky130_fd_sc_hd__dfxtp_1 _14887_ (.D(_02881_),
    .Q(\r1.regblock[26][4] ),
    .CLK(_01856_));
 sky130_fd_sc_hd__dfxtp_1 _14888_ (.D(_02882_),
    .Q(\r1.regblock[26][5] ),
    .CLK(_01857_));
 sky130_fd_sc_hd__dfxtp_1 _14889_ (.D(_02883_),
    .Q(\r1.regblock[26][6] ),
    .CLK(_01858_));
 sky130_fd_sc_hd__dfxtp_1 _14890_ (.D(_02884_),
    .Q(\r1.regblock[26][7] ),
    .CLK(_01859_));
 sky130_fd_sc_hd__dfxtp_1 _14891_ (.D(_02885_),
    .Q(\r1.regblock[26][8] ),
    .CLK(_01860_));
 sky130_fd_sc_hd__dfxtp_1 _14892_ (.D(_02886_),
    .Q(\r1.regblock[26][9] ),
    .CLK(_01861_));
 sky130_fd_sc_hd__dfxtp_1 _14893_ (.D(_02887_),
    .Q(\r1.regblock[26][10] ),
    .CLK(_01862_));
 sky130_fd_sc_hd__dfxtp_1 _14894_ (.D(_02888_),
    .Q(\r1.regblock[26][11] ),
    .CLK(_01863_));
 sky130_fd_sc_hd__dfxtp_1 _14895_ (.D(_02889_),
    .Q(\r1.regblock[26][12] ),
    .CLK(_01864_));
 sky130_fd_sc_hd__dfxtp_1 _14896_ (.D(_02890_),
    .Q(\r1.regblock[26][13] ),
    .CLK(_01865_));
 sky130_fd_sc_hd__dfxtp_1 _14897_ (.D(_02891_),
    .Q(\r1.regblock[26][14] ),
    .CLK(_01866_));
 sky130_fd_sc_hd__dfxtp_1 _14898_ (.D(_02892_),
    .Q(\r1.regblock[26][15] ),
    .CLK(_01867_));
 sky130_fd_sc_hd__dfxtp_1 _14899_ (.D(_02893_),
    .Q(\r1.regblock[26][16] ),
    .CLK(_01868_));
 sky130_fd_sc_hd__dfxtp_1 _14900_ (.D(_02894_),
    .Q(\r1.regblock[26][17] ),
    .CLK(_01869_));
 sky130_fd_sc_hd__dfxtp_1 _14901_ (.D(_02895_),
    .Q(\r1.regblock[26][18] ),
    .CLK(_01870_));
 sky130_fd_sc_hd__dfxtp_1 _14902_ (.D(_02896_),
    .Q(\r1.regblock[26][19] ),
    .CLK(_01871_));
 sky130_fd_sc_hd__dfxtp_1 _14903_ (.D(_02897_),
    .Q(\r1.regblock[26][20] ),
    .CLK(_01872_));
 sky130_fd_sc_hd__dfxtp_1 _14904_ (.D(_02898_),
    .Q(\r1.regblock[26][21] ),
    .CLK(_01873_));
 sky130_fd_sc_hd__dfxtp_1 _14905_ (.D(_02899_),
    .Q(\r1.regblock[26][22] ),
    .CLK(_01874_));
 sky130_fd_sc_hd__dfxtp_1 _14906_ (.D(_02900_),
    .Q(\r1.regblock[26][23] ),
    .CLK(_01875_));
 sky130_fd_sc_hd__dfxtp_1 _14907_ (.D(_02901_),
    .Q(\r1.regblock[26][24] ),
    .CLK(_01876_));
 sky130_fd_sc_hd__dfxtp_1 _14908_ (.D(_02902_),
    .Q(\r1.regblock[26][25] ),
    .CLK(_01877_));
 sky130_fd_sc_hd__dfxtp_1 _14909_ (.D(_02903_),
    .Q(\r1.regblock[26][26] ),
    .CLK(_01878_));
 sky130_fd_sc_hd__dfxtp_1 _14910_ (.D(_02904_),
    .Q(\r1.regblock[26][27] ),
    .CLK(_01879_));
 sky130_fd_sc_hd__dfxtp_1 _14911_ (.D(_02905_),
    .Q(\r1.regblock[26][28] ),
    .CLK(_01880_));
 sky130_fd_sc_hd__dfxtp_1 _14912_ (.D(_02906_),
    .Q(\r1.regblock[26][29] ),
    .CLK(_01881_));
 sky130_fd_sc_hd__dfxtp_1 _14913_ (.D(_02907_),
    .Q(\r1.regblock[26][30] ),
    .CLK(_01882_));
 sky130_fd_sc_hd__dfxtp_1 _14914_ (.D(_02908_),
    .Q(\r1.regblock[26][31] ),
    .CLK(_01883_));
 sky130_fd_sc_hd__dfxtp_1 _14915_ (.D(_02909_),
    .Q(\r1.regblock[27][0] ),
    .CLK(_01884_));
 sky130_fd_sc_hd__dfxtp_1 _14916_ (.D(_02910_),
    .Q(\r1.regblock[27][1] ),
    .CLK(_01885_));
 sky130_fd_sc_hd__dfxtp_1 _14917_ (.D(_02911_),
    .Q(\r1.regblock[27][2] ),
    .CLK(_01886_));
 sky130_fd_sc_hd__dfxtp_1 _14918_ (.D(_02912_),
    .Q(\r1.regblock[27][3] ),
    .CLK(_01887_));
 sky130_fd_sc_hd__dfxtp_1 _14919_ (.D(_02913_),
    .Q(\r1.regblock[27][4] ),
    .CLK(_01888_));
 sky130_fd_sc_hd__dfxtp_1 _14920_ (.D(_02914_),
    .Q(\r1.regblock[27][5] ),
    .CLK(_01889_));
 sky130_fd_sc_hd__dfxtp_1 _14921_ (.D(_02915_),
    .Q(\r1.regblock[27][6] ),
    .CLK(_01890_));
 sky130_fd_sc_hd__dfxtp_1 _14922_ (.D(_02916_),
    .Q(\r1.regblock[27][7] ),
    .CLK(_01891_));
 sky130_fd_sc_hd__dfxtp_1 _14923_ (.D(_02917_),
    .Q(\r1.regblock[27][8] ),
    .CLK(_01892_));
 sky130_fd_sc_hd__dfxtp_1 _14924_ (.D(_02918_),
    .Q(\r1.regblock[27][9] ),
    .CLK(_01893_));
 sky130_fd_sc_hd__dfxtp_1 _14925_ (.D(_02919_),
    .Q(\r1.regblock[27][10] ),
    .CLK(_01894_));
 sky130_fd_sc_hd__dfxtp_1 _14926_ (.D(_02920_),
    .Q(\r1.regblock[27][11] ),
    .CLK(_01895_));
 sky130_fd_sc_hd__dfxtp_1 _14927_ (.D(_02921_),
    .Q(\r1.regblock[27][12] ),
    .CLK(_01896_));
 sky130_fd_sc_hd__dfxtp_1 _14928_ (.D(_02922_),
    .Q(\r1.regblock[27][13] ),
    .CLK(_01897_));
 sky130_fd_sc_hd__dfxtp_1 _14929_ (.D(_02923_),
    .Q(\r1.regblock[27][14] ),
    .CLK(_01898_));
 sky130_fd_sc_hd__dfxtp_1 _14930_ (.D(_02924_),
    .Q(\r1.regblock[27][15] ),
    .CLK(_01899_));
 sky130_fd_sc_hd__dfxtp_1 _14931_ (.D(_02925_),
    .Q(\r1.regblock[27][16] ),
    .CLK(_01900_));
 sky130_fd_sc_hd__dfxtp_1 _14932_ (.D(_02926_),
    .Q(\r1.regblock[27][17] ),
    .CLK(_01901_));
 sky130_fd_sc_hd__dfxtp_1 _14933_ (.D(_02927_),
    .Q(\r1.regblock[27][18] ),
    .CLK(_01902_));
 sky130_fd_sc_hd__dfxtp_1 _14934_ (.D(_02928_),
    .Q(\r1.regblock[27][19] ),
    .CLK(_01903_));
 sky130_fd_sc_hd__dfxtp_1 _14935_ (.D(_02929_),
    .Q(\r1.regblock[27][20] ),
    .CLK(_01904_));
 sky130_fd_sc_hd__dfxtp_1 _14936_ (.D(_02930_),
    .Q(\r1.regblock[27][21] ),
    .CLK(_01905_));
 sky130_fd_sc_hd__dfxtp_1 _14937_ (.D(_02931_),
    .Q(\r1.regblock[27][22] ),
    .CLK(_01906_));
 sky130_fd_sc_hd__dfxtp_1 _14938_ (.D(_02932_),
    .Q(\r1.regblock[27][23] ),
    .CLK(_01907_));
 sky130_fd_sc_hd__dfxtp_1 _14939_ (.D(_02933_),
    .Q(\r1.regblock[27][24] ),
    .CLK(_01908_));
 sky130_fd_sc_hd__dfxtp_1 _14940_ (.D(_02934_),
    .Q(\r1.regblock[27][25] ),
    .CLK(_01909_));
 sky130_fd_sc_hd__dfxtp_1 _14941_ (.D(_02935_),
    .Q(\r1.regblock[27][26] ),
    .CLK(_01910_));
 sky130_fd_sc_hd__dfxtp_1 _14942_ (.D(_02936_),
    .Q(\r1.regblock[27][27] ),
    .CLK(_01911_));
 sky130_fd_sc_hd__dfxtp_1 _14943_ (.D(_02937_),
    .Q(\r1.regblock[27][28] ),
    .CLK(_01912_));
 sky130_fd_sc_hd__dfxtp_1 _14944_ (.D(_02938_),
    .Q(\r1.regblock[27][29] ),
    .CLK(_01913_));
 sky130_fd_sc_hd__dfxtp_1 _14945_ (.D(_02939_),
    .Q(\r1.regblock[27][30] ),
    .CLK(_01914_));
 sky130_fd_sc_hd__dfxtp_1 _14946_ (.D(_02940_),
    .Q(\r1.regblock[27][31] ),
    .CLK(_01915_));
 sky130_fd_sc_hd__dfxtp_1 _14947_ (.D(_02941_),
    .Q(\r1.regblock[28][0] ),
    .CLK(_01916_));
 sky130_fd_sc_hd__dfxtp_1 _14948_ (.D(_02942_),
    .Q(\r1.regblock[28][1] ),
    .CLK(_01917_));
 sky130_fd_sc_hd__dfxtp_1 _14949_ (.D(_02943_),
    .Q(\r1.regblock[28][2] ),
    .CLK(_01918_));
 sky130_fd_sc_hd__dfxtp_1 _14950_ (.D(_02944_),
    .Q(\r1.regblock[28][3] ),
    .CLK(_01919_));
 sky130_fd_sc_hd__dfxtp_1 _14951_ (.D(_02945_),
    .Q(\r1.regblock[28][4] ),
    .CLK(_01920_));
 sky130_fd_sc_hd__dfxtp_1 _14952_ (.D(_02946_),
    .Q(\r1.regblock[28][5] ),
    .CLK(_01921_));
 sky130_fd_sc_hd__dfxtp_1 _14953_ (.D(_02947_),
    .Q(\r1.regblock[28][6] ),
    .CLK(_01922_));
 sky130_fd_sc_hd__dfxtp_1 _14954_ (.D(_02948_),
    .Q(\r1.regblock[28][7] ),
    .CLK(_01923_));
 sky130_fd_sc_hd__dfxtp_1 _14955_ (.D(_02949_),
    .Q(\r1.regblock[28][8] ),
    .CLK(_01924_));
 sky130_fd_sc_hd__dfxtp_1 _14956_ (.D(_02950_),
    .Q(\r1.regblock[28][9] ),
    .CLK(_01925_));
 sky130_fd_sc_hd__dfxtp_1 _14957_ (.D(_02951_),
    .Q(\r1.regblock[28][10] ),
    .CLK(_01926_));
 sky130_fd_sc_hd__dfxtp_1 _14958_ (.D(_02952_),
    .Q(\r1.regblock[28][11] ),
    .CLK(_01927_));
 sky130_fd_sc_hd__dfxtp_1 _14959_ (.D(_02953_),
    .Q(\r1.regblock[28][12] ),
    .CLK(_01928_));
 sky130_fd_sc_hd__dfxtp_1 _14960_ (.D(_02954_),
    .Q(\r1.regblock[28][13] ),
    .CLK(_01929_));
 sky130_fd_sc_hd__dfxtp_1 _14961_ (.D(_02955_),
    .Q(\r1.regblock[28][14] ),
    .CLK(_01930_));
 sky130_fd_sc_hd__dfxtp_1 _14962_ (.D(_02956_),
    .Q(\r1.regblock[28][15] ),
    .CLK(_01931_));
 sky130_fd_sc_hd__dfxtp_1 _14963_ (.D(_02957_),
    .Q(\r1.regblock[28][16] ),
    .CLK(_01932_));
 sky130_fd_sc_hd__dfxtp_1 _14964_ (.D(_02958_),
    .Q(\r1.regblock[28][17] ),
    .CLK(_01933_));
 sky130_fd_sc_hd__dfxtp_1 _14965_ (.D(_02959_),
    .Q(\r1.regblock[28][18] ),
    .CLK(_01934_));
 sky130_fd_sc_hd__dfxtp_1 _14966_ (.D(_02960_),
    .Q(\r1.regblock[28][19] ),
    .CLK(_01935_));
 sky130_fd_sc_hd__dfxtp_1 _14967_ (.D(_02961_),
    .Q(\r1.regblock[28][20] ),
    .CLK(_01936_));
 sky130_fd_sc_hd__dfxtp_1 _14968_ (.D(_02962_),
    .Q(\r1.regblock[28][21] ),
    .CLK(_01937_));
 sky130_fd_sc_hd__dfxtp_1 _14969_ (.D(_02963_),
    .Q(\r1.regblock[28][22] ),
    .CLK(_01938_));
 sky130_fd_sc_hd__dfxtp_1 _14970_ (.D(_02964_),
    .Q(\r1.regblock[28][23] ),
    .CLK(_01939_));
 sky130_fd_sc_hd__dfxtp_1 _14971_ (.D(_02965_),
    .Q(\r1.regblock[28][24] ),
    .CLK(_01940_));
 sky130_fd_sc_hd__dfxtp_1 _14972_ (.D(_02966_),
    .Q(\r1.regblock[28][25] ),
    .CLK(_01941_));
 sky130_fd_sc_hd__dfxtp_1 _14973_ (.D(_02967_),
    .Q(\r1.regblock[28][26] ),
    .CLK(_01942_));
 sky130_fd_sc_hd__dfxtp_1 _14974_ (.D(_02968_),
    .Q(\r1.regblock[28][27] ),
    .CLK(_01943_));
 sky130_fd_sc_hd__dfxtp_1 _14975_ (.D(_02969_),
    .Q(\r1.regblock[28][28] ),
    .CLK(_01944_));
 sky130_fd_sc_hd__dfxtp_1 _14976_ (.D(_02970_),
    .Q(\r1.regblock[28][29] ),
    .CLK(_01945_));
 sky130_fd_sc_hd__dfxtp_1 _14977_ (.D(_02971_),
    .Q(\r1.regblock[28][30] ),
    .CLK(_01946_));
 sky130_fd_sc_hd__dfxtp_1 _14978_ (.D(_02972_),
    .Q(\r1.regblock[28][31] ),
    .CLK(_01947_));
 sky130_fd_sc_hd__dfxtp_1 _14979_ (.D(_02973_),
    .Q(\r1.regblock[2][0] ),
    .CLK(_01948_));
 sky130_fd_sc_hd__dfxtp_1 _14980_ (.D(_02974_),
    .Q(\r1.regblock[2][1] ),
    .CLK(_01949_));
 sky130_fd_sc_hd__dfxtp_1 _14981_ (.D(_02975_),
    .Q(\r1.regblock[2][2] ),
    .CLK(_01950_));
 sky130_fd_sc_hd__dfxtp_1 _14982_ (.D(_02976_),
    .Q(\r1.regblock[2][3] ),
    .CLK(_01951_));
 sky130_fd_sc_hd__dfxtp_1 _14983_ (.D(_02977_),
    .Q(\r1.regblock[2][4] ),
    .CLK(_01952_));
 sky130_fd_sc_hd__dfxtp_1 _14984_ (.D(_02978_),
    .Q(\r1.regblock[2][5] ),
    .CLK(_01953_));
 sky130_fd_sc_hd__dfxtp_1 _14985_ (.D(_02979_),
    .Q(\r1.regblock[2][6] ),
    .CLK(_01954_));
 sky130_fd_sc_hd__dfxtp_1 _14986_ (.D(_02980_),
    .Q(\r1.regblock[2][7] ),
    .CLK(_01955_));
 sky130_fd_sc_hd__dfxtp_1 _14987_ (.D(_02981_),
    .Q(\r1.regblock[2][8] ),
    .CLK(_01956_));
 sky130_fd_sc_hd__dfxtp_1 _14988_ (.D(_02982_),
    .Q(\r1.regblock[2][9] ),
    .CLK(_01957_));
 sky130_fd_sc_hd__dfxtp_1 _14989_ (.D(_02983_),
    .Q(\r1.regblock[2][10] ),
    .CLK(_01958_));
 sky130_fd_sc_hd__dfxtp_1 _14990_ (.D(_02984_),
    .Q(\r1.regblock[2][11] ),
    .CLK(_01959_));
 sky130_fd_sc_hd__dfxtp_1 _14991_ (.D(_02985_),
    .Q(\r1.regblock[2][12] ),
    .CLK(_01960_));
 sky130_fd_sc_hd__dfxtp_1 _14992_ (.D(_02986_),
    .Q(\r1.regblock[2][13] ),
    .CLK(_01961_));
 sky130_fd_sc_hd__dfxtp_1 _14993_ (.D(_02987_),
    .Q(\r1.regblock[2][14] ),
    .CLK(_01962_));
 sky130_fd_sc_hd__dfxtp_1 _14994_ (.D(_02988_),
    .Q(\r1.regblock[2][15] ),
    .CLK(_01963_));
 sky130_fd_sc_hd__dfxtp_1 _14995_ (.D(_02989_),
    .Q(\r1.regblock[2][16] ),
    .CLK(_01964_));
 sky130_fd_sc_hd__dfxtp_1 _14996_ (.D(_02990_),
    .Q(\r1.regblock[2][17] ),
    .CLK(_01965_));
 sky130_fd_sc_hd__dfxtp_1 _14997_ (.D(_02991_),
    .Q(\r1.regblock[2][18] ),
    .CLK(_01966_));
 sky130_fd_sc_hd__dfxtp_1 _14998_ (.D(_02992_),
    .Q(\r1.regblock[2][19] ),
    .CLK(_01967_));
 sky130_fd_sc_hd__dfxtp_1 _14999_ (.D(_02993_),
    .Q(\r1.regblock[2][20] ),
    .CLK(_01968_));
 sky130_fd_sc_hd__dfxtp_1 _15000_ (.D(_02994_),
    .Q(\r1.regblock[2][21] ),
    .CLK(_01969_));
 sky130_fd_sc_hd__dfxtp_1 _15001_ (.D(_02995_),
    .Q(\r1.regblock[2][22] ),
    .CLK(_01970_));
 sky130_fd_sc_hd__dfxtp_1 _15002_ (.D(_02996_),
    .Q(\r1.regblock[2][23] ),
    .CLK(_01971_));
 sky130_fd_sc_hd__dfxtp_1 _15003_ (.D(_02997_),
    .Q(\r1.regblock[2][24] ),
    .CLK(_01972_));
 sky130_fd_sc_hd__dfxtp_1 _15004_ (.D(_02998_),
    .Q(\r1.regblock[2][25] ),
    .CLK(_01973_));
 sky130_fd_sc_hd__dfxtp_1 _15005_ (.D(_02999_),
    .Q(\r1.regblock[2][26] ),
    .CLK(_01974_));
 sky130_fd_sc_hd__dfxtp_1 _15006_ (.D(_03000_),
    .Q(\r1.regblock[2][27] ),
    .CLK(_01975_));
 sky130_fd_sc_hd__dfxtp_1 _15007_ (.D(_03001_),
    .Q(\r1.regblock[2][28] ),
    .CLK(_01976_));
 sky130_fd_sc_hd__dfxtp_1 _15008_ (.D(_03002_),
    .Q(\r1.regblock[2][29] ),
    .CLK(_01977_));
 sky130_fd_sc_hd__dfxtp_1 _15009_ (.D(_03003_),
    .Q(\r1.regblock[2][30] ),
    .CLK(_01978_));
 sky130_fd_sc_hd__dfxtp_1 _15010_ (.D(_03004_),
    .Q(\r1.regblock[2][31] ),
    .CLK(_01979_));
 sky130_fd_sc_hd__dfxtp_1 _15011_ (.D(_03005_),
    .Q(\r1.regblock[30][0] ),
    .CLK(_01980_));
 sky130_fd_sc_hd__dfxtp_1 _15012_ (.D(_03006_),
    .Q(\r1.regblock[30][1] ),
    .CLK(_01981_));
 sky130_fd_sc_hd__dfxtp_1 _15013_ (.D(_03007_),
    .Q(\r1.regblock[30][2] ),
    .CLK(_01982_));
 sky130_fd_sc_hd__dfxtp_1 _15014_ (.D(_03008_),
    .Q(\r1.regblock[30][3] ),
    .CLK(_01983_));
 sky130_fd_sc_hd__dfxtp_1 _15015_ (.D(_03009_),
    .Q(\r1.regblock[30][4] ),
    .CLK(_01984_));
 sky130_fd_sc_hd__dfxtp_1 _15016_ (.D(_03010_),
    .Q(\r1.regblock[30][5] ),
    .CLK(_01985_));
 sky130_fd_sc_hd__dfxtp_1 _15017_ (.D(_03011_),
    .Q(\r1.regblock[30][6] ),
    .CLK(_01986_));
 sky130_fd_sc_hd__dfxtp_1 _15018_ (.D(_03012_),
    .Q(\r1.regblock[30][7] ),
    .CLK(_01987_));
 sky130_fd_sc_hd__dfxtp_1 _15019_ (.D(_03013_),
    .Q(\r1.regblock[30][8] ),
    .CLK(_01988_));
 sky130_fd_sc_hd__dfxtp_1 _15020_ (.D(_03014_),
    .Q(\r1.regblock[30][9] ),
    .CLK(_01989_));
 sky130_fd_sc_hd__dfxtp_1 _15021_ (.D(_03015_),
    .Q(\r1.regblock[30][10] ),
    .CLK(_01990_));
 sky130_fd_sc_hd__dfxtp_1 _15022_ (.D(_03016_),
    .Q(\r1.regblock[30][11] ),
    .CLK(_01991_));
 sky130_fd_sc_hd__dfxtp_1 _15023_ (.D(_03017_),
    .Q(\r1.regblock[30][12] ),
    .CLK(_01992_));
 sky130_fd_sc_hd__dfxtp_1 _15024_ (.D(_03018_),
    .Q(\r1.regblock[30][13] ),
    .CLK(_01993_));
 sky130_fd_sc_hd__dfxtp_1 _15025_ (.D(_03019_),
    .Q(\r1.regblock[30][14] ),
    .CLK(_01994_));
 sky130_fd_sc_hd__dfxtp_1 _15026_ (.D(_03020_),
    .Q(\r1.regblock[30][15] ),
    .CLK(_01995_));
 sky130_fd_sc_hd__dfxtp_1 _15027_ (.D(_03021_),
    .Q(\r1.regblock[30][16] ),
    .CLK(_01996_));
 sky130_fd_sc_hd__dfxtp_1 _15028_ (.D(_03022_),
    .Q(\r1.regblock[30][17] ),
    .CLK(_01997_));
 sky130_fd_sc_hd__dfxtp_1 _15029_ (.D(_03023_),
    .Q(\r1.regblock[30][18] ),
    .CLK(_01998_));
 sky130_fd_sc_hd__dfxtp_1 _15030_ (.D(_03024_),
    .Q(\r1.regblock[30][19] ),
    .CLK(_01999_));
 sky130_fd_sc_hd__dfxtp_1 _15031_ (.D(_03025_),
    .Q(\r1.regblock[30][20] ),
    .CLK(_02000_));
 sky130_fd_sc_hd__dfxtp_1 _15032_ (.D(_03026_),
    .Q(\r1.regblock[30][21] ),
    .CLK(_02001_));
 sky130_fd_sc_hd__dfxtp_1 _15033_ (.D(_03027_),
    .Q(\r1.regblock[30][22] ),
    .CLK(_02002_));
 sky130_fd_sc_hd__dfxtp_1 _15034_ (.D(_03028_),
    .Q(\r1.regblock[30][23] ),
    .CLK(_02003_));
 sky130_fd_sc_hd__dfxtp_1 _15035_ (.D(_03029_),
    .Q(\r1.regblock[30][24] ),
    .CLK(_02004_));
 sky130_fd_sc_hd__dfxtp_1 _15036_ (.D(_03030_),
    .Q(\r1.regblock[30][25] ),
    .CLK(_02005_));
 sky130_fd_sc_hd__dfxtp_1 _15037_ (.D(_03031_),
    .Q(\r1.regblock[30][26] ),
    .CLK(_02006_));
 sky130_fd_sc_hd__dfxtp_1 _15038_ (.D(_03032_),
    .Q(\r1.regblock[30][27] ),
    .CLK(_02007_));
 sky130_fd_sc_hd__dfxtp_1 _15039_ (.D(_03033_),
    .Q(\r1.regblock[30][28] ),
    .CLK(_02008_));
 sky130_fd_sc_hd__dfxtp_1 _15040_ (.D(_03034_),
    .Q(\r1.regblock[30][29] ),
    .CLK(_02009_));
 sky130_fd_sc_hd__dfxtp_1 _15041_ (.D(_03035_),
    .Q(\r1.regblock[30][30] ),
    .CLK(_02010_));
 sky130_fd_sc_hd__dfxtp_1 _15042_ (.D(_03036_),
    .Q(\r1.regblock[30][31] ),
    .CLK(_02011_));
 sky130_fd_sc_hd__dfxtp_1 _15043_ (.D(_03037_),
    .Q(\r1.regblock[29][0] ),
    .CLK(_02012_));
 sky130_fd_sc_hd__dfxtp_1 _15044_ (.D(_03038_),
    .Q(\r1.regblock[29][1] ),
    .CLK(_02013_));
 sky130_fd_sc_hd__dfxtp_1 _15045_ (.D(_03039_),
    .Q(\r1.regblock[29][2] ),
    .CLK(_02014_));
 sky130_fd_sc_hd__dfxtp_1 _15046_ (.D(_03040_),
    .Q(\r1.regblock[29][3] ),
    .CLK(_02015_));
 sky130_fd_sc_hd__dfxtp_1 _15047_ (.D(_03041_),
    .Q(\r1.regblock[29][4] ),
    .CLK(_02016_));
 sky130_fd_sc_hd__dfxtp_1 _15048_ (.D(_03042_),
    .Q(\r1.regblock[29][5] ),
    .CLK(_02017_));
 sky130_fd_sc_hd__dfxtp_1 _15049_ (.D(_03043_),
    .Q(\r1.regblock[29][6] ),
    .CLK(_02018_));
 sky130_fd_sc_hd__dfxtp_1 _15050_ (.D(_03044_),
    .Q(\r1.regblock[29][7] ),
    .CLK(_02019_));
 sky130_fd_sc_hd__dfxtp_1 _15051_ (.D(_03045_),
    .Q(\r1.regblock[29][8] ),
    .CLK(_02020_));
 sky130_fd_sc_hd__dfxtp_1 _15052_ (.D(_03046_),
    .Q(\r1.regblock[29][9] ),
    .CLK(_02021_));
 sky130_fd_sc_hd__dfxtp_1 _15053_ (.D(_03047_),
    .Q(\r1.regblock[29][10] ),
    .CLK(_02022_));
 sky130_fd_sc_hd__dfxtp_1 _15054_ (.D(_03048_),
    .Q(\r1.regblock[29][11] ),
    .CLK(_02023_));
 sky130_fd_sc_hd__dfxtp_1 _15055_ (.D(_03049_),
    .Q(\r1.regblock[29][12] ),
    .CLK(_02024_));
 sky130_fd_sc_hd__dfxtp_1 _15056_ (.D(_03050_),
    .Q(\r1.regblock[29][13] ),
    .CLK(_02025_));
 sky130_fd_sc_hd__dfxtp_1 _15057_ (.D(_03051_),
    .Q(\r1.regblock[29][14] ),
    .CLK(_02026_));
 sky130_fd_sc_hd__dfxtp_1 _15058_ (.D(_03052_),
    .Q(\r1.regblock[29][15] ),
    .CLK(_02027_));
 sky130_fd_sc_hd__dfxtp_1 _15059_ (.D(_03053_),
    .Q(\r1.regblock[29][16] ),
    .CLK(_02028_));
 sky130_fd_sc_hd__dfxtp_1 _15060_ (.D(_03054_),
    .Q(\r1.regblock[29][17] ),
    .CLK(_02029_));
 sky130_fd_sc_hd__dfxtp_1 _15061_ (.D(_03055_),
    .Q(\r1.regblock[29][18] ),
    .CLK(_02030_));
 sky130_fd_sc_hd__dfxtp_1 _15062_ (.D(_03056_),
    .Q(\r1.regblock[29][19] ),
    .CLK(_02031_));
 sky130_fd_sc_hd__dfxtp_1 _15063_ (.D(_03057_),
    .Q(\r1.regblock[29][20] ),
    .CLK(_02032_));
 sky130_fd_sc_hd__dfxtp_1 _15064_ (.D(_03058_),
    .Q(\r1.regblock[29][21] ),
    .CLK(_02033_));
 sky130_fd_sc_hd__dfxtp_1 _15065_ (.D(_03059_),
    .Q(\r1.regblock[29][22] ),
    .CLK(_02034_));
 sky130_fd_sc_hd__dfxtp_1 _15066_ (.D(_03060_),
    .Q(\r1.regblock[29][23] ),
    .CLK(_02035_));
 sky130_fd_sc_hd__dfxtp_1 _15067_ (.D(_03061_),
    .Q(\r1.regblock[29][24] ),
    .CLK(_02036_));
 sky130_fd_sc_hd__dfxtp_1 _15068_ (.D(_03062_),
    .Q(\r1.regblock[29][25] ),
    .CLK(_02037_));
 sky130_fd_sc_hd__dfxtp_1 _15069_ (.D(_03063_),
    .Q(\r1.regblock[29][26] ),
    .CLK(_02038_));
 sky130_fd_sc_hd__dfxtp_1 _15070_ (.D(_03064_),
    .Q(\r1.regblock[29][27] ),
    .CLK(_02039_));
 sky130_fd_sc_hd__dfxtp_1 _15071_ (.D(_03065_),
    .Q(\r1.regblock[29][28] ),
    .CLK(_02040_));
 sky130_fd_sc_hd__dfxtp_1 _15072_ (.D(_03066_),
    .Q(\r1.regblock[29][29] ),
    .CLK(_02041_));
 sky130_fd_sc_hd__dfxtp_1 _15073_ (.D(_03067_),
    .Q(\r1.regblock[29][30] ),
    .CLK(_02042_));
 sky130_fd_sc_hd__dfxtp_1 _15074_ (.D(_03068_),
    .Q(\r1.regblock[29][31] ),
    .CLK(_02043_));
 sky130_fd_sc_hd__dfxtp_1 _15075_ (.D(_03069_),
    .Q(\r1.regblock[31][0] ),
    .CLK(_02044_));
 sky130_fd_sc_hd__dfxtp_1 _15076_ (.D(_03070_),
    .Q(\r1.regblock[31][1] ),
    .CLK(_02045_));
 sky130_fd_sc_hd__dfxtp_1 _15077_ (.D(_03071_),
    .Q(\r1.regblock[31][2] ),
    .CLK(_02046_));
 sky130_fd_sc_hd__dfxtp_1 _15078_ (.D(_03072_),
    .Q(\r1.regblock[31][3] ),
    .CLK(_02047_));
 sky130_fd_sc_hd__dfxtp_1 _15079_ (.D(_03073_),
    .Q(\r1.regblock[31][4] ),
    .CLK(_02048_));
 sky130_fd_sc_hd__dfxtp_1 _15080_ (.D(_03074_),
    .Q(\r1.regblock[31][5] ),
    .CLK(_02049_));
 sky130_fd_sc_hd__dfxtp_1 _15081_ (.D(_03075_),
    .Q(\r1.regblock[31][6] ),
    .CLK(_02050_));
 sky130_fd_sc_hd__dfxtp_1 _15082_ (.D(_03076_),
    .Q(\r1.regblock[31][7] ),
    .CLK(_02051_));
 sky130_fd_sc_hd__dfxtp_1 _15083_ (.D(_03077_),
    .Q(\r1.regblock[31][8] ),
    .CLK(_02052_));
 sky130_fd_sc_hd__dfxtp_1 _15084_ (.D(_03078_),
    .Q(\r1.regblock[31][9] ),
    .CLK(_02053_));
 sky130_fd_sc_hd__dfxtp_1 _15085_ (.D(_03079_),
    .Q(\r1.regblock[31][10] ),
    .CLK(_02054_));
 sky130_fd_sc_hd__dfxtp_1 _15086_ (.D(_03080_),
    .Q(\r1.regblock[31][11] ),
    .CLK(_02055_));
 sky130_fd_sc_hd__dfxtp_1 _15087_ (.D(_03081_),
    .Q(\r1.regblock[31][12] ),
    .CLK(_02056_));
 sky130_fd_sc_hd__dfxtp_1 _15088_ (.D(_03082_),
    .Q(\r1.regblock[31][13] ),
    .CLK(_02057_));
 sky130_fd_sc_hd__dfxtp_1 _15089_ (.D(_03083_),
    .Q(\r1.regblock[31][14] ),
    .CLK(_02058_));
 sky130_fd_sc_hd__dfxtp_1 _15090_ (.D(_03084_),
    .Q(\r1.regblock[31][15] ),
    .CLK(_02059_));
 sky130_fd_sc_hd__dfxtp_1 _15091_ (.D(_03085_),
    .Q(\r1.regblock[31][16] ),
    .CLK(_02060_));
 sky130_fd_sc_hd__dfxtp_1 _15092_ (.D(_03086_),
    .Q(\r1.regblock[31][17] ),
    .CLK(_02061_));
 sky130_fd_sc_hd__dfxtp_1 _15093_ (.D(_03087_),
    .Q(\r1.regblock[31][18] ),
    .CLK(_02062_));
 sky130_fd_sc_hd__dfxtp_1 _15094_ (.D(_03088_),
    .Q(\r1.regblock[31][19] ),
    .CLK(_02063_));
 sky130_fd_sc_hd__dfxtp_1 _15095_ (.D(_03089_),
    .Q(\r1.regblock[31][20] ),
    .CLK(_02064_));
 sky130_fd_sc_hd__dfxtp_1 _15096_ (.D(_03090_),
    .Q(\r1.regblock[31][21] ),
    .CLK(_02065_));
 sky130_fd_sc_hd__dfxtp_1 _15097_ (.D(_03091_),
    .Q(\r1.regblock[31][22] ),
    .CLK(_02066_));
 sky130_fd_sc_hd__dfxtp_1 _15098_ (.D(_03092_),
    .Q(\r1.regblock[31][23] ),
    .CLK(_02067_));
 sky130_fd_sc_hd__dfxtp_1 _15099_ (.D(_03093_),
    .Q(\r1.regblock[31][24] ),
    .CLK(_02068_));
 sky130_fd_sc_hd__dfxtp_1 _15100_ (.D(_03094_),
    .Q(\r1.regblock[31][25] ),
    .CLK(_02069_));
 sky130_fd_sc_hd__dfxtp_1 _15101_ (.D(_03095_),
    .Q(\r1.regblock[31][26] ),
    .CLK(_02070_));
 sky130_fd_sc_hd__dfxtp_1 _15102_ (.D(_03096_),
    .Q(\r1.regblock[31][27] ),
    .CLK(_02071_));
 sky130_fd_sc_hd__dfxtp_1 _15103_ (.D(_03097_),
    .Q(\r1.regblock[31][28] ),
    .CLK(_02072_));
 sky130_fd_sc_hd__dfxtp_1 _15104_ (.D(_03098_),
    .Q(\r1.regblock[31][29] ),
    .CLK(_02073_));
 sky130_fd_sc_hd__dfxtp_1 _15105_ (.D(_03099_),
    .Q(\r1.regblock[31][30] ),
    .CLK(_02074_));
 sky130_fd_sc_hd__dfxtp_1 _15106_ (.D(_03100_),
    .Q(\r1.regblock[31][31] ),
    .CLK(_02075_));
 sky130_fd_sc_hd__dfxtp_1 _15107_ (.D(_03101_),
    .Q(\r1.regblock[12][0] ),
    .CLK(_02076_));
 sky130_fd_sc_hd__dfxtp_1 _15108_ (.D(_03102_),
    .Q(\r1.regblock[12][1] ),
    .CLK(_02077_));
 sky130_fd_sc_hd__dfxtp_1 _15109_ (.D(_03103_),
    .Q(\r1.regblock[12][2] ),
    .CLK(_02078_));
 sky130_fd_sc_hd__dfxtp_1 _15110_ (.D(_03104_),
    .Q(\r1.regblock[12][3] ),
    .CLK(_02079_));
 sky130_fd_sc_hd__dfxtp_1 _15111_ (.D(_03105_),
    .Q(\r1.regblock[12][4] ),
    .CLK(_02080_));
 sky130_fd_sc_hd__dfxtp_1 _15112_ (.D(_03106_),
    .Q(\r1.regblock[12][5] ),
    .CLK(_02081_));
 sky130_fd_sc_hd__dfxtp_1 _15113_ (.D(_03107_),
    .Q(\r1.regblock[12][6] ),
    .CLK(_02082_));
 sky130_fd_sc_hd__dfxtp_1 _15114_ (.D(_03108_),
    .Q(\r1.regblock[12][7] ),
    .CLK(_02083_));
 sky130_fd_sc_hd__dfxtp_1 _15115_ (.D(_03109_),
    .Q(\r1.regblock[12][8] ),
    .CLK(_02084_));
 sky130_fd_sc_hd__dfxtp_1 _15116_ (.D(_03110_),
    .Q(\r1.regblock[12][9] ),
    .CLK(_02085_));
 sky130_fd_sc_hd__dfxtp_1 _15117_ (.D(_03111_),
    .Q(\r1.regblock[12][10] ),
    .CLK(_02086_));
 sky130_fd_sc_hd__dfxtp_1 _15118_ (.D(_03112_),
    .Q(\r1.regblock[12][11] ),
    .CLK(_02087_));
 sky130_fd_sc_hd__dfxtp_1 _15119_ (.D(_03113_),
    .Q(\r1.regblock[12][12] ),
    .CLK(_02088_));
 sky130_fd_sc_hd__dfxtp_1 _15120_ (.D(_03114_),
    .Q(\r1.regblock[12][13] ),
    .CLK(_02089_));
 sky130_fd_sc_hd__dfxtp_1 _15121_ (.D(_03115_),
    .Q(\r1.regblock[12][14] ),
    .CLK(_02090_));
 sky130_fd_sc_hd__dfxtp_1 _15122_ (.D(_03116_),
    .Q(\r1.regblock[12][15] ),
    .CLK(_02091_));
 sky130_fd_sc_hd__dfxtp_1 _15123_ (.D(_03117_),
    .Q(\r1.regblock[12][16] ),
    .CLK(_02092_));
 sky130_fd_sc_hd__dfxtp_1 _15124_ (.D(_03118_),
    .Q(\r1.regblock[12][17] ),
    .CLK(_02093_));
 sky130_fd_sc_hd__dfxtp_1 _15125_ (.D(_03119_),
    .Q(\r1.regblock[12][18] ),
    .CLK(_02094_));
 sky130_fd_sc_hd__dfxtp_1 _15126_ (.D(_03120_),
    .Q(\r1.regblock[12][19] ),
    .CLK(_02095_));
 sky130_fd_sc_hd__dfxtp_1 _15127_ (.D(_03121_),
    .Q(\r1.regblock[12][20] ),
    .CLK(_02096_));
 sky130_fd_sc_hd__dfxtp_1 _15128_ (.D(_03122_),
    .Q(\r1.regblock[12][21] ),
    .CLK(_02097_));
 sky130_fd_sc_hd__dfxtp_1 _15129_ (.D(_03123_),
    .Q(\r1.regblock[12][22] ),
    .CLK(_02098_));
 sky130_fd_sc_hd__dfxtp_1 _15130_ (.D(_03124_),
    .Q(\r1.regblock[12][23] ),
    .CLK(_02099_));
 sky130_fd_sc_hd__dfxtp_1 _15131_ (.D(_03125_),
    .Q(\r1.regblock[12][24] ),
    .CLK(_02100_));
 sky130_fd_sc_hd__dfxtp_1 _15132_ (.D(_03126_),
    .Q(\r1.regblock[12][25] ),
    .CLK(_02101_));
 sky130_fd_sc_hd__dfxtp_1 _15133_ (.D(_03127_),
    .Q(\r1.regblock[12][26] ),
    .CLK(_02102_));
 sky130_fd_sc_hd__dfxtp_1 _15134_ (.D(_03128_),
    .Q(\r1.regblock[12][27] ),
    .CLK(_02103_));
 sky130_fd_sc_hd__dfxtp_1 _15135_ (.D(_03129_),
    .Q(\r1.regblock[12][28] ),
    .CLK(_02104_));
 sky130_fd_sc_hd__dfxtp_1 _15136_ (.D(_03130_),
    .Q(\r1.regblock[12][29] ),
    .CLK(_02105_));
 sky130_fd_sc_hd__dfxtp_1 _15137_ (.D(_03131_),
    .Q(\r1.regblock[12][30] ),
    .CLK(_02106_));
 sky130_fd_sc_hd__dfxtp_1 _15138_ (.D(_03132_),
    .Q(\r1.regblock[12][31] ),
    .CLK(_02107_));
 sky130_fd_sc_hd__dfxtp_1 _15139_ (.D(_03133_),
    .Q(\r1.regblock[9][0] ),
    .CLK(_02108_));
 sky130_fd_sc_hd__dfxtp_1 _15140_ (.D(_03134_),
    .Q(\r1.regblock[9][1] ),
    .CLK(_02109_));
 sky130_fd_sc_hd__dfxtp_1 _15141_ (.D(_03135_),
    .Q(\r1.regblock[9][2] ),
    .CLK(_02110_));
 sky130_fd_sc_hd__dfxtp_1 _15142_ (.D(_03136_),
    .Q(\r1.regblock[9][3] ),
    .CLK(_02111_));
 sky130_fd_sc_hd__dfxtp_1 _15143_ (.D(_03137_),
    .Q(\r1.regblock[9][4] ),
    .CLK(_02112_));
 sky130_fd_sc_hd__dfxtp_1 _15144_ (.D(_03138_),
    .Q(\r1.regblock[9][5] ),
    .CLK(_02113_));
 sky130_fd_sc_hd__dfxtp_1 _15145_ (.D(_03139_),
    .Q(\r1.regblock[9][6] ),
    .CLK(_02114_));
 sky130_fd_sc_hd__dfxtp_1 _15146_ (.D(_03140_),
    .Q(\r1.regblock[9][7] ),
    .CLK(_02115_));
 sky130_fd_sc_hd__dfxtp_1 _15147_ (.D(_03141_),
    .Q(\r1.regblock[9][8] ),
    .CLK(_02116_));
 sky130_fd_sc_hd__dfxtp_1 _15148_ (.D(_03142_),
    .Q(\r1.regblock[9][9] ),
    .CLK(_02117_));
 sky130_fd_sc_hd__dfxtp_1 _15149_ (.D(_03143_),
    .Q(\r1.regblock[9][10] ),
    .CLK(_02118_));
 sky130_fd_sc_hd__dfxtp_1 _15150_ (.D(_03144_),
    .Q(\r1.regblock[9][11] ),
    .CLK(_02119_));
 sky130_fd_sc_hd__dfxtp_1 _15151_ (.D(_03145_),
    .Q(\r1.regblock[9][12] ),
    .CLK(_02120_));
 sky130_fd_sc_hd__dfxtp_1 _15152_ (.D(_03146_),
    .Q(\r1.regblock[9][13] ),
    .CLK(_02121_));
 sky130_fd_sc_hd__dfxtp_1 _15153_ (.D(_03147_),
    .Q(\r1.regblock[9][14] ),
    .CLK(_02122_));
 sky130_fd_sc_hd__dfxtp_1 _15154_ (.D(_03148_),
    .Q(\r1.regblock[9][15] ),
    .CLK(_02123_));
 sky130_fd_sc_hd__dfxtp_1 _15155_ (.D(_03149_),
    .Q(\r1.regblock[9][16] ),
    .CLK(_02124_));
 sky130_fd_sc_hd__dfxtp_1 _15156_ (.D(_03150_),
    .Q(\r1.regblock[9][17] ),
    .CLK(_02125_));
 sky130_fd_sc_hd__dfxtp_1 _15157_ (.D(_03151_),
    .Q(\r1.regblock[9][18] ),
    .CLK(_02126_));
 sky130_fd_sc_hd__dfxtp_1 _15158_ (.D(_03152_),
    .Q(\r1.regblock[9][19] ),
    .CLK(_02127_));
 sky130_fd_sc_hd__dfxtp_1 _15159_ (.D(_03153_),
    .Q(\r1.regblock[9][20] ),
    .CLK(_02128_));
 sky130_fd_sc_hd__dfxtp_1 _15160_ (.D(_03154_),
    .Q(\r1.regblock[9][21] ),
    .CLK(_02129_));
 sky130_fd_sc_hd__dfxtp_1 _15161_ (.D(_03155_),
    .Q(\r1.regblock[9][22] ),
    .CLK(_02130_));
 sky130_fd_sc_hd__dfxtp_1 _15162_ (.D(_03156_),
    .Q(\r1.regblock[9][23] ),
    .CLK(_02131_));
 sky130_fd_sc_hd__dfxtp_1 _15163_ (.D(_03157_),
    .Q(\r1.regblock[9][24] ),
    .CLK(_02132_));
 sky130_fd_sc_hd__dfxtp_1 _15164_ (.D(_03158_),
    .Q(\r1.regblock[9][25] ),
    .CLK(_02133_));
 sky130_fd_sc_hd__dfxtp_1 _15165_ (.D(_03159_),
    .Q(\r1.regblock[9][26] ),
    .CLK(_02134_));
 sky130_fd_sc_hd__dfxtp_1 _15166_ (.D(_03160_),
    .Q(\r1.regblock[9][27] ),
    .CLK(_02135_));
 sky130_fd_sc_hd__dfxtp_1 _15167_ (.D(_03161_),
    .Q(\r1.regblock[9][28] ),
    .CLK(_02136_));
 sky130_fd_sc_hd__dfxtp_1 _15168_ (.D(_03162_),
    .Q(\r1.regblock[9][29] ),
    .CLK(_02137_));
 sky130_fd_sc_hd__dfxtp_1 _15169_ (.D(_03163_),
    .Q(\r1.regblock[9][30] ),
    .CLK(_02138_));
 sky130_fd_sc_hd__dfxtp_1 _15170_ (.D(_03164_),
    .Q(\r1.regblock[9][31] ),
    .CLK(_02139_));
 sky130_fd_sc_hd__dfxtp_1 _15171_ (.D(_03165_),
    .Q(\r1.regblock[8][0] ),
    .CLK(_02140_));
 sky130_fd_sc_hd__dfxtp_1 _15172_ (.D(_03166_),
    .Q(\r1.regblock[8][1] ),
    .CLK(_02141_));
 sky130_fd_sc_hd__dfxtp_1 _15173_ (.D(_03167_),
    .Q(\r1.regblock[8][2] ),
    .CLK(_02142_));
 sky130_fd_sc_hd__dfxtp_1 _15174_ (.D(_03168_),
    .Q(\r1.regblock[8][3] ),
    .CLK(_02143_));
 sky130_fd_sc_hd__dfxtp_1 _15175_ (.D(_03169_),
    .Q(\r1.regblock[8][4] ),
    .CLK(_02144_));
 sky130_fd_sc_hd__dfxtp_1 _15176_ (.D(_03170_),
    .Q(\r1.regblock[8][5] ),
    .CLK(_02145_));
 sky130_fd_sc_hd__dfxtp_1 _15177_ (.D(_03171_),
    .Q(\r1.regblock[8][6] ),
    .CLK(_02146_));
 sky130_fd_sc_hd__dfxtp_1 _15178_ (.D(_03172_),
    .Q(\r1.regblock[8][7] ),
    .CLK(_02147_));
 sky130_fd_sc_hd__dfxtp_1 _15179_ (.D(_03173_),
    .Q(\r1.regblock[8][8] ),
    .CLK(_02148_));
 sky130_fd_sc_hd__dfxtp_1 _15180_ (.D(_03174_),
    .Q(\r1.regblock[8][9] ),
    .CLK(_02149_));
 sky130_fd_sc_hd__dfxtp_1 _15181_ (.D(_03175_),
    .Q(\r1.regblock[8][10] ),
    .CLK(_02150_));
 sky130_fd_sc_hd__dfxtp_1 _15182_ (.D(_03176_),
    .Q(\r1.regblock[8][11] ),
    .CLK(_02151_));
 sky130_fd_sc_hd__dfxtp_1 _15183_ (.D(_03177_),
    .Q(\r1.regblock[8][12] ),
    .CLK(_02152_));
 sky130_fd_sc_hd__dfxtp_1 _15184_ (.D(_03178_),
    .Q(\r1.regblock[8][13] ),
    .CLK(_02153_));
 sky130_fd_sc_hd__dfxtp_1 _15185_ (.D(_03179_),
    .Q(\r1.regblock[8][14] ),
    .CLK(_02154_));
 sky130_fd_sc_hd__dfxtp_1 _15186_ (.D(_03180_),
    .Q(\r1.regblock[8][15] ),
    .CLK(_02155_));
 sky130_fd_sc_hd__dfxtp_1 _15187_ (.D(_03181_),
    .Q(\r1.regblock[8][16] ),
    .CLK(_02156_));
 sky130_fd_sc_hd__dfxtp_1 _15188_ (.D(_03182_),
    .Q(\r1.regblock[8][17] ),
    .CLK(_02157_));
 sky130_fd_sc_hd__dfxtp_1 _15189_ (.D(_03183_),
    .Q(\r1.regblock[8][18] ),
    .CLK(_02158_));
 sky130_fd_sc_hd__dfxtp_1 _15190_ (.D(_03184_),
    .Q(\r1.regblock[8][19] ),
    .CLK(_02159_));
 sky130_fd_sc_hd__dfxtp_1 _15191_ (.D(_03185_),
    .Q(\r1.regblock[8][20] ),
    .CLK(_02160_));
 sky130_fd_sc_hd__dfxtp_1 _15192_ (.D(_03186_),
    .Q(\r1.regblock[8][21] ),
    .CLK(_02161_));
 sky130_fd_sc_hd__dfxtp_1 _15193_ (.D(_03187_),
    .Q(\r1.regblock[8][22] ),
    .CLK(_02162_));
 sky130_fd_sc_hd__dfxtp_1 _15194_ (.D(_03188_),
    .Q(\r1.regblock[8][23] ),
    .CLK(_02163_));
 sky130_fd_sc_hd__dfxtp_1 _15195_ (.D(_03189_),
    .Q(\r1.regblock[8][24] ),
    .CLK(_02164_));
 sky130_fd_sc_hd__dfxtp_1 _15196_ (.D(_03190_),
    .Q(\r1.regblock[8][25] ),
    .CLK(_02165_));
 sky130_fd_sc_hd__dfxtp_1 _15197_ (.D(_03191_),
    .Q(\r1.regblock[8][26] ),
    .CLK(_02166_));
 sky130_fd_sc_hd__dfxtp_1 _15198_ (.D(_03192_),
    .Q(\r1.regblock[8][27] ),
    .CLK(_02167_));
 sky130_fd_sc_hd__dfxtp_1 _15199_ (.D(_03193_),
    .Q(\r1.regblock[8][28] ),
    .CLK(_02168_));
 sky130_fd_sc_hd__dfxtp_1 _15200_ (.D(_03194_),
    .Q(\r1.regblock[8][29] ),
    .CLK(_02169_));
 sky130_fd_sc_hd__dfxtp_1 _15201_ (.D(_03195_),
    .Q(\r1.regblock[8][30] ),
    .CLK(_02170_));
 sky130_fd_sc_hd__dfxtp_1 _15202_ (.D(_03196_),
    .Q(\r1.regblock[8][31] ),
    .CLK(_02171_));
 sky130_fd_sc_hd__dfxtp_1 _15203_ (.D(_03197_),
    .Q(\r1.regblock[0][0] ),
    .CLK(_02172_));
 sky130_fd_sc_hd__dfxtp_1 _15204_ (.D(_03198_),
    .Q(\r1.regblock[0][1] ),
    .CLK(_02173_));
 sky130_fd_sc_hd__dfxtp_1 _15205_ (.D(_03199_),
    .Q(\r1.regblock[0][2] ),
    .CLK(_02174_));
 sky130_fd_sc_hd__dfxtp_1 _15206_ (.D(_03200_),
    .Q(\r1.regblock[0][3] ),
    .CLK(_02175_));
 sky130_fd_sc_hd__dfxtp_1 _15207_ (.D(_03201_),
    .Q(\r1.regblock[0][4] ),
    .CLK(_02176_));
 sky130_fd_sc_hd__dfxtp_1 _15208_ (.D(_03202_),
    .Q(\r1.regblock[0][5] ),
    .CLK(_02177_));
 sky130_fd_sc_hd__dfxtp_1 _15209_ (.D(_03203_),
    .Q(\r1.regblock[0][6] ),
    .CLK(_02178_));
 sky130_fd_sc_hd__dfxtp_1 _15210_ (.D(_03204_),
    .Q(\r1.regblock[0][7] ),
    .CLK(_02179_));
 sky130_fd_sc_hd__dfxtp_1 _15211_ (.D(_03205_),
    .Q(\r1.regblock[0][8] ),
    .CLK(_02180_));
 sky130_fd_sc_hd__dfxtp_1 _15212_ (.D(_03206_),
    .Q(\r1.regblock[0][9] ),
    .CLK(_02181_));
 sky130_fd_sc_hd__dfxtp_1 _15213_ (.D(_03207_),
    .Q(\r1.regblock[0][10] ),
    .CLK(_02182_));
 sky130_fd_sc_hd__dfxtp_1 _15214_ (.D(_03208_),
    .Q(\r1.regblock[0][11] ),
    .CLK(_02183_));
 sky130_fd_sc_hd__dfxtp_1 _15215_ (.D(_03209_),
    .Q(\r1.regblock[0][12] ),
    .CLK(_02184_));
 sky130_fd_sc_hd__dfxtp_1 _15216_ (.D(_03210_),
    .Q(\r1.regblock[0][13] ),
    .CLK(_02185_));
 sky130_fd_sc_hd__dfxtp_1 _15217_ (.D(_03211_),
    .Q(\r1.regblock[0][14] ),
    .CLK(_02186_));
 sky130_fd_sc_hd__dfxtp_1 _15218_ (.D(_03212_),
    .Q(\r1.regblock[0][15] ),
    .CLK(_02187_));
 sky130_fd_sc_hd__dfxtp_1 _15219_ (.D(_03213_),
    .Q(\r1.regblock[0][16] ),
    .CLK(_02188_));
 sky130_fd_sc_hd__dfxtp_1 _15220_ (.D(_03214_),
    .Q(\r1.regblock[0][17] ),
    .CLK(_02189_));
 sky130_fd_sc_hd__dfxtp_1 _15221_ (.D(_03215_),
    .Q(\r1.regblock[0][18] ),
    .CLK(_02190_));
 sky130_fd_sc_hd__dfxtp_1 _15222_ (.D(_03216_),
    .Q(\r1.regblock[0][19] ),
    .CLK(_02191_));
 sky130_fd_sc_hd__dfxtp_1 _15223_ (.D(_03217_),
    .Q(\r1.regblock[0][20] ),
    .CLK(_02192_));
 sky130_fd_sc_hd__dfxtp_1 _15224_ (.D(_03218_),
    .Q(\r1.regblock[0][21] ),
    .CLK(_02193_));
 sky130_fd_sc_hd__dfxtp_1 _15225_ (.D(_03219_),
    .Q(\r1.regblock[0][22] ),
    .CLK(_02194_));
 sky130_fd_sc_hd__dfxtp_1 _15226_ (.D(_03220_),
    .Q(\r1.regblock[0][23] ),
    .CLK(_02195_));
 sky130_fd_sc_hd__dfxtp_1 _15227_ (.D(_03221_),
    .Q(\r1.regblock[0][24] ),
    .CLK(_02196_));
 sky130_fd_sc_hd__dfxtp_1 _15228_ (.D(_03222_),
    .Q(\r1.regblock[0][25] ),
    .CLK(_02197_));
 sky130_fd_sc_hd__dfxtp_1 _15229_ (.D(_03223_),
    .Q(\r1.regblock[0][26] ),
    .CLK(_02198_));
 sky130_fd_sc_hd__dfxtp_1 _15230_ (.D(_03224_),
    .Q(\r1.regblock[0][27] ),
    .CLK(_02199_));
 sky130_fd_sc_hd__dfxtp_1 _15231_ (.D(_03225_),
    .Q(\r1.regblock[0][28] ),
    .CLK(_02200_));
 sky130_fd_sc_hd__dfxtp_1 _15232_ (.D(_03226_),
    .Q(\r1.regblock[0][29] ),
    .CLK(_02201_));
 sky130_fd_sc_hd__dfxtp_1 _15233_ (.D(_03227_),
    .Q(\r1.regblock[0][30] ),
    .CLK(_02202_));
 sky130_fd_sc_hd__dfxtp_1 _15234_ (.D(_03228_),
    .Q(\r1.regblock[0][31] ),
    .CLK(_02203_));
 sky130_fd_sc_hd__dfxtp_1 _15235_ (.D(_03229_),
    .Q(\r1.regblock[5][0] ),
    .CLK(_02204_));
 sky130_fd_sc_hd__dfxtp_1 _15236_ (.D(_03230_),
    .Q(\r1.regblock[5][1] ),
    .CLK(_02205_));
 sky130_fd_sc_hd__dfxtp_1 _15237_ (.D(_03231_),
    .Q(\r1.regblock[5][2] ),
    .CLK(_02206_));
 sky130_fd_sc_hd__dfxtp_1 _15238_ (.D(_03232_),
    .Q(\r1.regblock[5][3] ),
    .CLK(_02207_));
 sky130_fd_sc_hd__dfxtp_1 _15239_ (.D(_03233_),
    .Q(\r1.regblock[5][4] ),
    .CLK(_02208_));
 sky130_fd_sc_hd__dfxtp_1 _15240_ (.D(_03234_),
    .Q(\r1.regblock[5][5] ),
    .CLK(_02209_));
 sky130_fd_sc_hd__dfxtp_1 _15241_ (.D(_03235_),
    .Q(\r1.regblock[5][6] ),
    .CLK(_02210_));
 sky130_fd_sc_hd__dfxtp_1 _15242_ (.D(_03236_),
    .Q(\r1.regblock[5][7] ),
    .CLK(_02211_));
 sky130_fd_sc_hd__dfxtp_1 _15243_ (.D(_03237_),
    .Q(\r1.regblock[5][8] ),
    .CLK(_02212_));
 sky130_fd_sc_hd__dfxtp_1 _15244_ (.D(_03238_),
    .Q(\r1.regblock[5][9] ),
    .CLK(_02213_));
 sky130_fd_sc_hd__dfxtp_1 _15245_ (.D(_03239_),
    .Q(\r1.regblock[5][10] ),
    .CLK(_02214_));
 sky130_fd_sc_hd__dfxtp_1 _15246_ (.D(_03240_),
    .Q(\r1.regblock[5][11] ),
    .CLK(_02215_));
 sky130_fd_sc_hd__dfxtp_1 _15247_ (.D(_03241_),
    .Q(\r1.regblock[5][12] ),
    .CLK(_02216_));
 sky130_fd_sc_hd__dfxtp_1 _15248_ (.D(_03242_),
    .Q(\r1.regblock[5][13] ),
    .CLK(_02217_));
 sky130_fd_sc_hd__dfxtp_1 _15249_ (.D(_03243_),
    .Q(\r1.regblock[5][14] ),
    .CLK(_02218_));
 sky130_fd_sc_hd__dfxtp_1 _15250_ (.D(_03244_),
    .Q(\r1.regblock[5][15] ),
    .CLK(_02219_));
 sky130_fd_sc_hd__dfxtp_1 _15251_ (.D(_03245_),
    .Q(\r1.regblock[5][16] ),
    .CLK(_02220_));
 sky130_fd_sc_hd__dfxtp_1 _15252_ (.D(_03246_),
    .Q(\r1.regblock[5][17] ),
    .CLK(_02221_));
 sky130_fd_sc_hd__dfxtp_1 _15253_ (.D(_03247_),
    .Q(\r1.regblock[5][18] ),
    .CLK(_02222_));
 sky130_fd_sc_hd__dfxtp_1 _15254_ (.D(_03248_),
    .Q(\r1.regblock[5][19] ),
    .CLK(_02223_));
 sky130_fd_sc_hd__dfxtp_1 _15255_ (.D(_03249_),
    .Q(\r1.regblock[5][20] ),
    .CLK(_02224_));
 sky130_fd_sc_hd__dfxtp_1 _15256_ (.D(_03250_),
    .Q(\r1.regblock[5][21] ),
    .CLK(_02225_));
 sky130_fd_sc_hd__dfxtp_1 _15257_ (.D(_03251_),
    .Q(\r1.regblock[5][22] ),
    .CLK(_02226_));
 sky130_fd_sc_hd__dfxtp_1 _15258_ (.D(_03252_),
    .Q(\r1.regblock[5][23] ),
    .CLK(_02227_));
 sky130_fd_sc_hd__dfxtp_1 _15259_ (.D(_03253_),
    .Q(\r1.regblock[5][24] ),
    .CLK(_02228_));
 sky130_fd_sc_hd__dfxtp_1 _15260_ (.D(_03254_),
    .Q(\r1.regblock[5][25] ),
    .CLK(_02229_));
 sky130_fd_sc_hd__dfxtp_1 _15261_ (.D(_03255_),
    .Q(\r1.regblock[5][26] ),
    .CLK(_02230_));
 sky130_fd_sc_hd__dfxtp_1 _15262_ (.D(_03256_),
    .Q(\r1.regblock[5][27] ),
    .CLK(_02231_));
 sky130_fd_sc_hd__dfxtp_1 _15263_ (.D(_03257_),
    .Q(\r1.regblock[5][28] ),
    .CLK(_02232_));
 sky130_fd_sc_hd__dfxtp_1 _15264_ (.D(_03258_),
    .Q(\r1.regblock[5][29] ),
    .CLK(_02233_));
 sky130_fd_sc_hd__dfxtp_1 _15265_ (.D(_03259_),
    .Q(\r1.regblock[5][30] ),
    .CLK(_02234_));
 sky130_fd_sc_hd__dfxtp_1 _15266_ (.D(_03260_),
    .Q(\r1.regblock[5][31] ),
    .CLK(_02235_));
 sky130_fd_sc_hd__dfxtp_1 _15267_ (.D(_03261_),
    .Q(\r1.regblock[15][0] ),
    .CLK(_02236_));
 sky130_fd_sc_hd__dfxtp_1 _15268_ (.D(_03262_),
    .Q(\r1.regblock[15][1] ),
    .CLK(_02237_));
 sky130_fd_sc_hd__dfxtp_1 _15269_ (.D(_03263_),
    .Q(\r1.regblock[15][2] ),
    .CLK(_02238_));
 sky130_fd_sc_hd__dfxtp_1 _15270_ (.D(_03264_),
    .Q(\r1.regblock[15][3] ),
    .CLK(_02239_));
 sky130_fd_sc_hd__dfxtp_1 _15271_ (.D(_03265_),
    .Q(\r1.regblock[15][4] ),
    .CLK(_02240_));
 sky130_fd_sc_hd__dfxtp_1 _15272_ (.D(_03266_),
    .Q(\r1.regblock[15][5] ),
    .CLK(_02241_));
 sky130_fd_sc_hd__dfxtp_1 _15273_ (.D(_03267_),
    .Q(\r1.regblock[15][6] ),
    .CLK(_02242_));
 sky130_fd_sc_hd__dfxtp_1 _15274_ (.D(_03268_),
    .Q(\r1.regblock[15][7] ),
    .CLK(_02243_));
 sky130_fd_sc_hd__dfxtp_1 _15275_ (.D(_03269_),
    .Q(\r1.regblock[15][8] ),
    .CLK(_02244_));
 sky130_fd_sc_hd__dfxtp_1 _15276_ (.D(_03270_),
    .Q(\r1.regblock[15][9] ),
    .CLK(_02245_));
 sky130_fd_sc_hd__dfxtp_1 _15277_ (.D(_03271_),
    .Q(\r1.regblock[15][10] ),
    .CLK(_02246_));
 sky130_fd_sc_hd__dfxtp_1 _15278_ (.D(_03272_),
    .Q(\r1.regblock[15][11] ),
    .CLK(_02247_));
 sky130_fd_sc_hd__dfxtp_1 _15279_ (.D(_03273_),
    .Q(\r1.regblock[15][12] ),
    .CLK(_02248_));
 sky130_fd_sc_hd__dfxtp_1 _15280_ (.D(_03274_),
    .Q(\r1.regblock[15][13] ),
    .CLK(_02249_));
 sky130_fd_sc_hd__dfxtp_1 _15281_ (.D(_03275_),
    .Q(\r1.regblock[15][14] ),
    .CLK(_02250_));
 sky130_fd_sc_hd__dfxtp_1 _15282_ (.D(_03276_),
    .Q(\r1.regblock[15][15] ),
    .CLK(_02251_));
 sky130_fd_sc_hd__dfxtp_1 _15283_ (.D(_03277_),
    .Q(\r1.regblock[15][16] ),
    .CLK(_02252_));
 sky130_fd_sc_hd__dfxtp_1 _15284_ (.D(_03278_),
    .Q(\r1.regblock[15][17] ),
    .CLK(_02253_));
 sky130_fd_sc_hd__dfxtp_1 _15285_ (.D(_03279_),
    .Q(\r1.regblock[15][18] ),
    .CLK(_02254_));
 sky130_fd_sc_hd__dfxtp_1 _15286_ (.D(_03280_),
    .Q(\r1.regblock[15][19] ),
    .CLK(_02255_));
 sky130_fd_sc_hd__dfxtp_1 _15287_ (.D(_03281_),
    .Q(\r1.regblock[15][20] ),
    .CLK(_02256_));
 sky130_fd_sc_hd__dfxtp_1 _15288_ (.D(_03282_),
    .Q(\r1.regblock[15][21] ),
    .CLK(_02257_));
 sky130_fd_sc_hd__dfxtp_1 _15289_ (.D(_03283_),
    .Q(\r1.regblock[15][22] ),
    .CLK(_02258_));
 sky130_fd_sc_hd__dfxtp_1 _15290_ (.D(_03284_),
    .Q(\r1.regblock[15][23] ),
    .CLK(_02259_));
 sky130_fd_sc_hd__dfxtp_1 _15291_ (.D(_03285_),
    .Q(\r1.regblock[15][24] ),
    .CLK(_02260_));
 sky130_fd_sc_hd__dfxtp_1 _15292_ (.D(_03286_),
    .Q(\r1.regblock[15][25] ),
    .CLK(_02261_));
 sky130_fd_sc_hd__dfxtp_1 _15293_ (.D(_03287_),
    .Q(\r1.regblock[15][26] ),
    .CLK(_02262_));
 sky130_fd_sc_hd__dfxtp_1 _15294_ (.D(_03288_),
    .Q(\r1.regblock[15][27] ),
    .CLK(_02263_));
 sky130_fd_sc_hd__dfxtp_1 _15295_ (.D(_03289_),
    .Q(\r1.regblock[15][28] ),
    .CLK(_02264_));
 sky130_fd_sc_hd__dfxtp_1 _15296_ (.D(_03290_),
    .Q(\r1.regblock[15][29] ),
    .CLK(_02265_));
 sky130_fd_sc_hd__dfxtp_1 _15297_ (.D(_03291_),
    .Q(\r1.regblock[15][30] ),
    .CLK(_02266_));
 sky130_fd_sc_hd__dfxtp_1 _15298_ (.D(_03292_),
    .Q(\r1.regblock[15][31] ),
    .CLK(_02267_));
 sky130_fd_sc_hd__dfxtp_1 _15299_ (.D(_03293_),
    .Q(\r1.regblock[14][0] ),
    .CLK(_02268_));
 sky130_fd_sc_hd__dfxtp_1 _15300_ (.D(_03294_),
    .Q(\r1.regblock[14][1] ),
    .CLK(_02269_));
 sky130_fd_sc_hd__dfxtp_1 _15301_ (.D(_03295_),
    .Q(\r1.regblock[14][2] ),
    .CLK(_02270_));
 sky130_fd_sc_hd__dfxtp_1 _15302_ (.D(_03296_),
    .Q(\r1.regblock[14][3] ),
    .CLK(_02271_));
 sky130_fd_sc_hd__dfxtp_1 _15303_ (.D(_03297_),
    .Q(\r1.regblock[14][4] ),
    .CLK(_02272_));
 sky130_fd_sc_hd__dfxtp_1 _15304_ (.D(_03298_),
    .Q(\r1.regblock[14][5] ),
    .CLK(_02273_));
 sky130_fd_sc_hd__dfxtp_1 _15305_ (.D(_03299_),
    .Q(\r1.regblock[14][6] ),
    .CLK(_02274_));
 sky130_fd_sc_hd__dfxtp_1 _15306_ (.D(_03300_),
    .Q(\r1.regblock[14][7] ),
    .CLK(_02275_));
 sky130_fd_sc_hd__dfxtp_1 _15307_ (.D(_03301_),
    .Q(\r1.regblock[14][8] ),
    .CLK(_02276_));
 sky130_fd_sc_hd__dfxtp_1 _15308_ (.D(_03302_),
    .Q(\r1.regblock[14][9] ),
    .CLK(_02277_));
 sky130_fd_sc_hd__dfxtp_1 _15309_ (.D(_03303_),
    .Q(\r1.regblock[14][10] ),
    .CLK(_02278_));
 sky130_fd_sc_hd__dfxtp_1 _15310_ (.D(_03304_),
    .Q(\r1.regblock[14][11] ),
    .CLK(_02279_));
 sky130_fd_sc_hd__dfxtp_1 _15311_ (.D(_03305_),
    .Q(\r1.regblock[14][12] ),
    .CLK(_02280_));
 sky130_fd_sc_hd__dfxtp_1 _15312_ (.D(_03306_),
    .Q(\r1.regblock[14][13] ),
    .CLK(_02281_));
 sky130_fd_sc_hd__dfxtp_1 _15313_ (.D(_03307_),
    .Q(\r1.regblock[14][14] ),
    .CLK(_02282_));
 sky130_fd_sc_hd__dfxtp_1 _15314_ (.D(_03308_),
    .Q(\r1.regblock[14][15] ),
    .CLK(_02283_));
 sky130_fd_sc_hd__dfxtp_1 _15315_ (.D(_03309_),
    .Q(\r1.regblock[14][16] ),
    .CLK(_02284_));
 sky130_fd_sc_hd__dfxtp_1 _15316_ (.D(_03310_),
    .Q(\r1.regblock[14][17] ),
    .CLK(_02285_));
 sky130_fd_sc_hd__dfxtp_1 _15317_ (.D(_03311_),
    .Q(\r1.regblock[14][18] ),
    .CLK(_02286_));
 sky130_fd_sc_hd__dfxtp_1 _15318_ (.D(_03312_),
    .Q(\r1.regblock[14][19] ),
    .CLK(_02287_));
 sky130_fd_sc_hd__dfxtp_1 _15319_ (.D(_03313_),
    .Q(\r1.regblock[14][20] ),
    .CLK(_02288_));
 sky130_fd_sc_hd__dfxtp_1 _15320_ (.D(_03314_),
    .Q(\r1.regblock[14][21] ),
    .CLK(_02289_));
 sky130_fd_sc_hd__dfxtp_1 _15321_ (.D(_03315_),
    .Q(\r1.regblock[14][22] ),
    .CLK(_02290_));
 sky130_fd_sc_hd__dfxtp_1 _15322_ (.D(_03316_),
    .Q(\r1.regblock[14][23] ),
    .CLK(_02291_));
 sky130_fd_sc_hd__dfxtp_1 _15323_ (.D(_03317_),
    .Q(\r1.regblock[14][24] ),
    .CLK(_02292_));
 sky130_fd_sc_hd__dfxtp_1 _15324_ (.D(_03318_),
    .Q(\r1.regblock[14][25] ),
    .CLK(_02293_));
 sky130_fd_sc_hd__dfxtp_1 _15325_ (.D(_03319_),
    .Q(\r1.regblock[14][26] ),
    .CLK(_02294_));
 sky130_fd_sc_hd__dfxtp_1 _15326_ (.D(_03320_),
    .Q(\r1.regblock[14][27] ),
    .CLK(_02295_));
 sky130_fd_sc_hd__dfxtp_1 _15327_ (.D(_03321_),
    .Q(\r1.regblock[14][28] ),
    .CLK(_02296_));
 sky130_fd_sc_hd__dfxtp_1 _15328_ (.D(_03322_),
    .Q(\r1.regblock[14][29] ),
    .CLK(_02297_));
 sky130_fd_sc_hd__dfxtp_1 _15329_ (.D(_03323_),
    .Q(\r1.regblock[14][30] ),
    .CLK(_02298_));
 sky130_fd_sc_hd__dfxtp_1 _15330_ (.D(_03324_),
    .Q(\r1.regblock[14][31] ),
    .CLK(_02299_));
 sky130_fd_sc_hd__dfxtp_1 _15331_ (.D(_03325_),
    .Q(\r1.regblock[13][0] ),
    .CLK(_02300_));
 sky130_fd_sc_hd__dfxtp_1 _15332_ (.D(_03326_),
    .Q(\r1.regblock[13][1] ),
    .CLK(_02301_));
 sky130_fd_sc_hd__dfxtp_1 _15333_ (.D(_03327_),
    .Q(\r1.regblock[13][2] ),
    .CLK(_02302_));
 sky130_fd_sc_hd__dfxtp_1 _15334_ (.D(_03328_),
    .Q(\r1.regblock[13][3] ),
    .CLK(_02303_));
 sky130_fd_sc_hd__dfxtp_1 _15335_ (.D(_03329_),
    .Q(\r1.regblock[13][4] ),
    .CLK(_02304_));
 sky130_fd_sc_hd__dfxtp_1 _15336_ (.D(_03330_),
    .Q(\r1.regblock[13][5] ),
    .CLK(_02305_));
 sky130_fd_sc_hd__dfxtp_1 _15337_ (.D(_03331_),
    .Q(\r1.regblock[13][6] ),
    .CLK(_02306_));
 sky130_fd_sc_hd__dfxtp_1 _15338_ (.D(_03332_),
    .Q(\r1.regblock[13][7] ),
    .CLK(_02307_));
 sky130_fd_sc_hd__dfxtp_1 _15339_ (.D(_03333_),
    .Q(\r1.regblock[13][8] ),
    .CLK(_02308_));
 sky130_fd_sc_hd__dfxtp_1 _15340_ (.D(_03334_),
    .Q(\r1.regblock[13][9] ),
    .CLK(_02309_));
 sky130_fd_sc_hd__dfxtp_1 _15341_ (.D(_03335_),
    .Q(\r1.regblock[13][10] ),
    .CLK(_02310_));
 sky130_fd_sc_hd__dfxtp_1 _15342_ (.D(_03336_),
    .Q(\r1.regblock[13][11] ),
    .CLK(_02311_));
 sky130_fd_sc_hd__dfxtp_1 _15343_ (.D(_03337_),
    .Q(\r1.regblock[13][12] ),
    .CLK(_02312_));
 sky130_fd_sc_hd__dfxtp_1 _15344_ (.D(_03338_),
    .Q(\r1.regblock[13][13] ),
    .CLK(_02313_));
 sky130_fd_sc_hd__dfxtp_1 _15345_ (.D(_03339_),
    .Q(\r1.regblock[13][14] ),
    .CLK(_02314_));
 sky130_fd_sc_hd__dfxtp_1 _15346_ (.D(_03340_),
    .Q(\r1.regblock[13][15] ),
    .CLK(_02315_));
 sky130_fd_sc_hd__dfxtp_1 _15347_ (.D(_03341_),
    .Q(\r1.regblock[13][16] ),
    .CLK(_02316_));
 sky130_fd_sc_hd__dfxtp_1 _15348_ (.D(_03342_),
    .Q(\r1.regblock[13][17] ),
    .CLK(_02317_));
 sky130_fd_sc_hd__dfxtp_1 _15349_ (.D(_03343_),
    .Q(\r1.regblock[13][18] ),
    .CLK(_02318_));
 sky130_fd_sc_hd__dfxtp_1 _15350_ (.D(_03344_),
    .Q(\r1.regblock[13][19] ),
    .CLK(_02319_));
 sky130_fd_sc_hd__dfxtp_1 _15351_ (.D(_03345_),
    .Q(\r1.regblock[13][20] ),
    .CLK(_02320_));
 sky130_fd_sc_hd__dfxtp_1 _15352_ (.D(_03346_),
    .Q(\r1.regblock[13][21] ),
    .CLK(_02321_));
 sky130_fd_sc_hd__dfxtp_1 _15353_ (.D(_03347_),
    .Q(\r1.regblock[13][22] ),
    .CLK(_02322_));
 sky130_fd_sc_hd__dfxtp_1 _15354_ (.D(_03348_),
    .Q(\r1.regblock[13][23] ),
    .CLK(_02323_));
 sky130_fd_sc_hd__dfxtp_1 _15355_ (.D(_03349_),
    .Q(\r1.regblock[13][24] ),
    .CLK(_02324_));
 sky130_fd_sc_hd__dfxtp_1 _15356_ (.D(_03350_),
    .Q(\r1.regblock[13][25] ),
    .CLK(_02325_));
 sky130_fd_sc_hd__dfxtp_1 _15357_ (.D(_03351_),
    .Q(\r1.regblock[13][26] ),
    .CLK(_02326_));
 sky130_fd_sc_hd__dfxtp_1 _15358_ (.D(_03352_),
    .Q(\r1.regblock[13][27] ),
    .CLK(_02327_));
 sky130_fd_sc_hd__dfxtp_1 _15359_ (.D(_03353_),
    .Q(\r1.regblock[13][28] ),
    .CLK(_02328_));
 sky130_fd_sc_hd__dfxtp_1 _15360_ (.D(_03354_),
    .Q(\r1.regblock[13][29] ),
    .CLK(_02329_));
 sky130_fd_sc_hd__dfxtp_1 _15361_ (.D(_03355_),
    .Q(\r1.regblock[13][30] ),
    .CLK(_02330_));
 sky130_fd_sc_hd__dfxtp_1 _15362_ (.D(_03356_),
    .Q(\r1.regblock[13][31] ),
    .CLK(_02331_));
 sky130_fd_sc_hd__dfxtp_1 _15363_ (.D(_03357_),
    .Q(\r1.regblock[19][0] ),
    .CLK(_02332_));
 sky130_fd_sc_hd__dfxtp_1 _15364_ (.D(_03358_),
    .Q(\r1.regblock[19][1] ),
    .CLK(_02333_));
 sky130_fd_sc_hd__dfxtp_1 _15365_ (.D(_03359_),
    .Q(\r1.regblock[19][2] ),
    .CLK(_02334_));
 sky130_fd_sc_hd__dfxtp_1 _15366_ (.D(_03360_),
    .Q(\r1.regblock[19][3] ),
    .CLK(_02335_));
 sky130_fd_sc_hd__dfxtp_1 _15367_ (.D(_03361_),
    .Q(\r1.regblock[19][4] ),
    .CLK(_02336_));
 sky130_fd_sc_hd__dfxtp_1 _15368_ (.D(_03362_),
    .Q(\r1.regblock[19][5] ),
    .CLK(_02337_));
 sky130_fd_sc_hd__dfxtp_1 _15369_ (.D(_03363_),
    .Q(\r1.regblock[19][6] ),
    .CLK(_02338_));
 sky130_fd_sc_hd__dfxtp_1 _15370_ (.D(_03364_),
    .Q(\r1.regblock[19][7] ),
    .CLK(_02339_));
 sky130_fd_sc_hd__dfxtp_1 _15371_ (.D(_03365_),
    .Q(\r1.regblock[19][8] ),
    .CLK(_02340_));
 sky130_fd_sc_hd__dfxtp_1 _15372_ (.D(_03366_),
    .Q(\r1.regblock[19][9] ),
    .CLK(_02341_));
 sky130_fd_sc_hd__dfxtp_1 _15373_ (.D(_03367_),
    .Q(\r1.regblock[19][10] ),
    .CLK(_02342_));
 sky130_fd_sc_hd__dfxtp_1 _15374_ (.D(_03368_),
    .Q(\r1.regblock[19][11] ),
    .CLK(_02343_));
 sky130_fd_sc_hd__dfxtp_1 _15375_ (.D(_03369_),
    .Q(\r1.regblock[19][12] ),
    .CLK(_02344_));
 sky130_fd_sc_hd__dfxtp_1 _15376_ (.D(_03370_),
    .Q(\r1.regblock[19][13] ),
    .CLK(_02345_));
 sky130_fd_sc_hd__dfxtp_1 _15377_ (.D(_03371_),
    .Q(\r1.regblock[19][14] ),
    .CLK(_02346_));
 sky130_fd_sc_hd__dfxtp_1 _15378_ (.D(_03372_),
    .Q(\r1.regblock[19][15] ),
    .CLK(_02347_));
 sky130_fd_sc_hd__dfxtp_1 _15379_ (.D(_03373_),
    .Q(\r1.regblock[19][16] ),
    .CLK(_02348_));
 sky130_fd_sc_hd__dfxtp_1 _15380_ (.D(_03374_),
    .Q(\r1.regblock[19][17] ),
    .CLK(_02349_));
 sky130_fd_sc_hd__dfxtp_1 _15381_ (.D(_03375_),
    .Q(\r1.regblock[19][18] ),
    .CLK(_02350_));
 sky130_fd_sc_hd__dfxtp_1 _15382_ (.D(_03376_),
    .Q(\r1.regblock[19][19] ),
    .CLK(_02351_));
 sky130_fd_sc_hd__dfxtp_1 _15383_ (.D(_03377_),
    .Q(\r1.regblock[19][20] ),
    .CLK(_02352_));
 sky130_fd_sc_hd__dfxtp_1 _15384_ (.D(_03378_),
    .Q(\r1.regblock[19][21] ),
    .CLK(_02353_));
 sky130_fd_sc_hd__dfxtp_1 _15385_ (.D(_03379_),
    .Q(\r1.regblock[19][22] ),
    .CLK(_02354_));
 sky130_fd_sc_hd__dfxtp_1 _15386_ (.D(_03380_),
    .Q(\r1.regblock[19][23] ),
    .CLK(_02355_));
 sky130_fd_sc_hd__dfxtp_1 _15387_ (.D(_03381_),
    .Q(\r1.regblock[19][24] ),
    .CLK(_02356_));
 sky130_fd_sc_hd__dfxtp_1 _15388_ (.D(_03382_),
    .Q(\r1.regblock[19][25] ),
    .CLK(_02357_));
 sky130_fd_sc_hd__dfxtp_1 _15389_ (.D(_03383_),
    .Q(\r1.regblock[19][26] ),
    .CLK(_02358_));
 sky130_fd_sc_hd__dfxtp_1 _15390_ (.D(_03384_),
    .Q(\r1.regblock[19][27] ),
    .CLK(_02359_));
 sky130_fd_sc_hd__dfxtp_1 _15391_ (.D(_03385_),
    .Q(\r1.regblock[19][28] ),
    .CLK(_02360_));
 sky130_fd_sc_hd__dfxtp_1 _15392_ (.D(_03386_),
    .Q(\r1.regblock[19][29] ),
    .CLK(_02361_));
 sky130_fd_sc_hd__dfxtp_1 _15393_ (.D(_03387_),
    .Q(\r1.regblock[19][30] ),
    .CLK(_02362_));
 sky130_fd_sc_hd__dfxtp_1 _15394_ (.D(_03388_),
    .Q(\r1.regblock[19][31] ),
    .CLK(_02363_));
 sky130_fd_sc_hd__dfxtp_1 _15395_ (.D(_03389_),
    .Q(\r1.regblock[3][0] ),
    .CLK(_02364_));
 sky130_fd_sc_hd__dfxtp_1 _15396_ (.D(_03390_),
    .Q(\r1.regblock[3][1] ),
    .CLK(_02365_));
 sky130_fd_sc_hd__dfxtp_1 _15397_ (.D(_03391_),
    .Q(\r1.regblock[3][2] ),
    .CLK(_02366_));
 sky130_fd_sc_hd__dfxtp_1 _15398_ (.D(_03392_),
    .Q(\r1.regblock[3][3] ),
    .CLK(_02367_));
 sky130_fd_sc_hd__dfxtp_1 _15399_ (.D(_03393_),
    .Q(\r1.regblock[3][4] ),
    .CLK(_02368_));
 sky130_fd_sc_hd__dfxtp_1 _15400_ (.D(_03394_),
    .Q(\r1.regblock[3][5] ),
    .CLK(_02369_));
 sky130_fd_sc_hd__dfxtp_1 _15401_ (.D(_03395_),
    .Q(\r1.regblock[3][6] ),
    .CLK(_02370_));
 sky130_fd_sc_hd__dfxtp_1 _15402_ (.D(_03396_),
    .Q(\r1.regblock[3][7] ),
    .CLK(_02371_));
 sky130_fd_sc_hd__dfxtp_1 _15403_ (.D(_03397_),
    .Q(\r1.regblock[3][8] ),
    .CLK(_02372_));
 sky130_fd_sc_hd__dfxtp_1 _15404_ (.D(_03398_),
    .Q(\r1.regblock[3][9] ),
    .CLK(_02373_));
 sky130_fd_sc_hd__dfxtp_1 _15405_ (.D(_03399_),
    .Q(\r1.regblock[3][10] ),
    .CLK(_02374_));
 sky130_fd_sc_hd__dfxtp_1 _15406_ (.D(_03400_),
    .Q(\r1.regblock[3][11] ),
    .CLK(_02375_));
 sky130_fd_sc_hd__dfxtp_1 _15407_ (.D(_03401_),
    .Q(\r1.regblock[3][12] ),
    .CLK(_02376_));
 sky130_fd_sc_hd__dfxtp_1 _15408_ (.D(_03402_),
    .Q(\r1.regblock[3][13] ),
    .CLK(_02377_));
 sky130_fd_sc_hd__dfxtp_1 _15409_ (.D(_03403_),
    .Q(\r1.regblock[3][14] ),
    .CLK(_02378_));
 sky130_fd_sc_hd__dfxtp_1 _15410_ (.D(_03404_),
    .Q(\r1.regblock[3][15] ),
    .CLK(_02379_));
 sky130_fd_sc_hd__dfxtp_1 _15411_ (.D(_03405_),
    .Q(\r1.regblock[3][16] ),
    .CLK(_02380_));
 sky130_fd_sc_hd__dfxtp_1 _15412_ (.D(_03406_),
    .Q(\r1.regblock[3][17] ),
    .CLK(_02381_));
 sky130_fd_sc_hd__dfxtp_1 _15413_ (.D(_03407_),
    .Q(\r1.regblock[3][18] ),
    .CLK(_02382_));
 sky130_fd_sc_hd__dfxtp_1 _15414_ (.D(_03408_),
    .Q(\r1.regblock[3][19] ),
    .CLK(_02383_));
 sky130_fd_sc_hd__dfxtp_1 _15415_ (.D(_03409_),
    .Q(\r1.regblock[3][20] ),
    .CLK(_02384_));
 sky130_fd_sc_hd__dfxtp_1 _15416_ (.D(_03410_),
    .Q(\r1.regblock[3][21] ),
    .CLK(_02385_));
 sky130_fd_sc_hd__dfxtp_1 _15417_ (.D(_03411_),
    .Q(\r1.regblock[3][22] ),
    .CLK(_02386_));
 sky130_fd_sc_hd__dfxtp_1 _15418_ (.D(_03412_),
    .Q(\r1.regblock[3][23] ),
    .CLK(_02387_));
 sky130_fd_sc_hd__dfxtp_1 _15419_ (.D(_03413_),
    .Q(\r1.regblock[3][24] ),
    .CLK(_02388_));
 sky130_fd_sc_hd__dfxtp_1 _15420_ (.D(_03414_),
    .Q(\r1.regblock[3][25] ),
    .CLK(_02389_));
 sky130_fd_sc_hd__dfxtp_1 _15421_ (.D(_03415_),
    .Q(\r1.regblock[3][26] ),
    .CLK(_02390_));
 sky130_fd_sc_hd__dfxtp_1 _15422_ (.D(_03416_),
    .Q(\r1.regblock[3][27] ),
    .CLK(_02391_));
 sky130_fd_sc_hd__dfxtp_1 _15423_ (.D(_03417_),
    .Q(\r1.regblock[3][28] ),
    .CLK(_02392_));
 sky130_fd_sc_hd__dfxtp_1 _15424_ (.D(_03418_),
    .Q(\r1.regblock[3][29] ),
    .CLK(_02393_));
 sky130_fd_sc_hd__dfxtp_1 _15425_ (.D(_03419_),
    .Q(\r1.regblock[3][30] ),
    .CLK(_02394_));
 sky130_fd_sc_hd__dfxtp_1 _15426_ (.D(_03420_),
    .Q(\r1.regblock[3][31] ),
    .CLK(_02395_));
 sky130_fd_sc_hd__dfxtp_4 _15427_ (.D(_03421_),
    .Q(data_address[0]),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_2 _15428_ (.D(_03422_),
    .Q(data_address[1]),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_4 _15429_ (.D(_03423_),
    .Q(data_address[2]),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_4 _15430_ (.D(_03424_),
    .Q(data_address[3]),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_4 _15431_ (.D(_03425_),
    .Q(data_address[4]),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _15432_ (.D(_03426_),
    .Q(data_address[5]),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_2 _15433_ (.D(_03427_),
    .Q(data_address[6]),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_4 _15434_ (.D(_03428_),
    .Q(data_address[7]),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_4 _15435_ (.D(_03429_),
    .Q(data_address[8]),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_2 _15436_ (.D(_03430_),
    .Q(data_address[9]),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_4 _15437_ (.D(_03431_),
    .Q(data_address[10]),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _15438_ (.D(_03432_),
    .Q(data_address[11]),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_4 _15439_ (.D(_03433_),
    .Q(data_address[12]),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 _15440_ (.D(_03434_),
    .Q(data_address[13]),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_4 _15441_ (.D(_03435_),
    .Q(data_address[14]),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _15442_ (.D(_03436_),
    .Q(data_address[15]),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_4 _15443_ (.D(_03437_),
    .Q(data_address[16]),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 _15444_ (.D(_03438_),
    .Q(data_address[17]),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_4 _15445_ (.D(_03439_),
    .Q(data_address[18]),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 _15446_ (.D(_03440_),
    .Q(data_address[19]),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_2 _15447_ (.D(_03441_),
    .Q(data_address[20]),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_2 _15448_ (.D(_03442_),
    .Q(data_address[21]),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_4 _15449_ (.D(_03443_),
    .Q(data_address[22]),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _15450_ (.D(_03444_),
    .Q(data_address[23]),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _15451_ (.D(_03445_),
    .Q(data_address[24]),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _15452_ (.D(_03446_),
    .Q(data_address[25]),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _15453_ (.D(_03447_),
    .Q(data_address[26]),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_4 _15454_ (.D(_03448_),
    .Q(data_address[27]),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_4 _15455_ (.D(_03449_),
    .Q(data_address[28]),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_4 _15456_ (.D(_03450_),
    .Q(data_address[29]),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _15457_ (.D(_03451_),
    .Q(data_address[30]),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _15458_ (.D(_03452_),
    .Q(data_address[31]),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 _15459_ (.D(_03453_),
    .Q(\c1.instruction3[0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _15460_ (.D(_03454_),
    .Q(\c1.instruction3[1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _15461_ (.D(_03455_),
    .Q(\c1.instruction3[2] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _15462_ (.D(_03456_),
    .Q(\c1.instruction3[3] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _15463_ (.D(_03457_),
    .Q(\c1.instruction3[4] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _15464_ (.D(_03458_),
    .Q(\c1.instruction3[5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _15465_ (.D(_03459_),
    .Q(\c1.instruction3[6] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _15466_ (.D(_03460_),
    .Q(\c1.instruction3[7] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 _15467_ (.D(_03461_),
    .Q(\c1.instruction3[8] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _15468_ (.D(_03462_),
    .Q(\c1.instruction3[9] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _15469_ (.D(_03463_),
    .Q(\c1.instruction3[10] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _15470_ (.D(_03464_),
    .Q(\c1.instruction3[11] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _15471_ (.D(_03465_),
    .Q(\c1.instruction3[12] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _15472_ (.D(_03466_),
    .Q(\c1.instruction3[13] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _15473_ (.D(_03467_),
    .Q(\c1.instruction3[14] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_2 _15474_ (.D(_03468_),
    .Q(wdata[0]),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_2 _15475_ (.D(_03469_),
    .Q(wdata[1]),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _15476_ (.D(_03470_),
    .Q(wdata[2]),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _15477_ (.D(_03471_),
    .Q(wdata[3]),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_4 _15478_ (.D(_03472_),
    .Q(wdata[4]),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_4 _15479_ (.D(_03473_),
    .Q(wdata[5]),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _15480_ (.D(_03474_),
    .Q(wdata[6]),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _15481_ (.D(_03475_),
    .Q(wdata[7]),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _15482_ (.D(_03476_),
    .Q(wdata[8]),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _15483_ (.D(_03477_),
    .Q(wdata[9]),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_4 _15484_ (.D(_03478_),
    .Q(wdata[10]),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_4 _15485_ (.D(_03479_),
    .Q(wdata[11]),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _15486_ (.D(_03480_),
    .Q(wdata[12]),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_4 _15487_ (.D(_03481_),
    .Q(wdata[13]),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_2 _15488_ (.D(_03482_),
    .Q(wdata[14]),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_2 _15489_ (.D(_03483_),
    .Q(wdata[15]),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_2 _15490_ (.D(_03484_),
    .Q(wdata[16]),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 _15491_ (.D(_03485_),
    .Q(wdata[17]),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 _15492_ (.D(_03486_),
    .Q(wdata[18]),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_4 _15493_ (.D(_03487_),
    .Q(wdata[19]),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_4 _15494_ (.D(_03488_),
    .Q(wdata[20]),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_2 _15495_ (.D(_03489_),
    .Q(wdata[21]),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_4 _15496_ (.D(_03490_),
    .Q(wdata[22]),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _15497_ (.D(_03491_),
    .Q(wdata[23]),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_4 _15498_ (.D(_03492_),
    .Q(wdata[24]),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 _15499_ (.D(_03493_),
    .Q(wdata[25]),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _15500_ (.D(_03494_),
    .Q(wdata[26]),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _15501_ (.D(_03495_),
    .Q(wdata[27]),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _15502_ (.D(_03496_),
    .Q(wdata[28]),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_4 _15503_ (.D(_03497_),
    .Q(wdata[29]),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _15504_ (.D(_03498_),
    .Q(wdata[30]),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_2 _15505_ (.D(_03499_),
    .Q(wdata[31]),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_4 _15506_ (.D(_03500_),
    .Q(\DEP_PLACE[3] ),
    .CLK(_02396_));
 sky130_fd_sc_hd__dfxtp_1 _15507_ (.D(_03501_),
    .Q(\c1.instruction2[0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _15508_ (.D(_03502_),
    .Q(\c1.instruction2[1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _15509_ (.D(_03503_),
    .Q(\c1.instruction2[2] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 _15510_ (.D(_03504_),
    .Q(\c1.instruction2[3] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _15511_ (.D(_03505_),
    .Q(\c1.instruction2[4] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _15512_ (.D(_03506_),
    .Q(\c1.instruction2[5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _15513_ (.D(_03507_),
    .Q(\c1.instruction2[6] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 _15514_ (.D(_03508_),
    .Q(\c1.instruction2[7] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 _15515_ (.D(_03509_),
    .Q(\c1.instruction2[8] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _15516_ (.D(_03510_),
    .Q(\c1.instruction2[9] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _15517_ (.D(_03511_),
    .Q(\c1.instruction2[10] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _15518_ (.D(_03512_),
    .Q(\c1.instruction2[11] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _15519_ (.D(_03513_),
    .Q(\c1.instruction2[12] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _15520_ (.D(_03514_),
    .Q(\c1.instruction2[13] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _15521_ (.D(_03515_),
    .Q(\c1.instruction2[14] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _15522_ (.D(_03516_),
    .Q(\c1.instruction2[25] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 _15523_ (.D(_03517_),
    .Q(\c1.instruction2[26] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 _15524_ (.D(_03518_),
    .Q(\c1.instruction2[27] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 _15525_ (.D(_03519_),
    .Q(\c1.instruction2[28] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 _15526_ (.D(_03520_),
    .Q(\c1.instruction2[29] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 _15527_ (.D(_03521_),
    .Q(\c1.instruction2[30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 _15528_ (.D(_03522_),
    .Q(\c1.instruction2[31] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _15529_ (.D(_03523_),
    .Q(\e1.alu1.a[0] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _15530_ (.D(_03524_),
    .Q(\e1.alu1.a[1] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15531_ (.D(_03525_),
    .Q(\e1.alu1.a[2] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15532_ (.D(_03526_),
    .Q(\e1.alu1.a[3] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15533_ (.D(_03527_),
    .Q(\e1.alu1.a[4] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15534_ (.D(_03528_),
    .Q(\e1.alu1.a[5] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _15535_ (.D(_03529_),
    .Q(\e1.alu1.a[6] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _15536_ (.D(_03530_),
    .Q(\e1.alu1.a[7] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15537_ (.D(_03531_),
    .Q(\e1.alu1.a[8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _15538_ (.D(_03532_),
    .Q(\e1.alu1.a[9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _15539_ (.D(_03533_),
    .Q(\e1.alu1.a[10] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _15540_ (.D(_03534_),
    .Q(\e1.alu1.a[11] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 _15541_ (.D(_03535_),
    .Q(\e1.alu1.a[12] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _15542_ (.D(_03536_),
    .Q(\e1.alu1.a[13] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _15543_ (.D(_03537_),
    .Q(\e1.alu1.a[14] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 _15544_ (.D(_03538_),
    .Q(\e1.alu1.a[15] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 _15545_ (.D(_03539_),
    .Q(\e1.alu1.a[16] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15546_ (.D(_03540_),
    .Q(\e1.alu1.a[17] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _15547_ (.D(_03541_),
    .Q(\e1.alu1.a[18] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _15548_ (.D(_03542_),
    .Q(\e1.alu1.a[19] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _15549_ (.D(_03543_),
    .Q(\e1.alu1.a[20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _15550_ (.D(_03544_),
    .Q(\e1.alu1.a[21] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _15551_ (.D(_03545_),
    .Q(\e1.alu1.a[22] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _15552_ (.D(_03546_),
    .Q(\e1.alu1.a[23] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _15553_ (.D(_03547_),
    .Q(\e1.alu1.a[24] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _15554_ (.D(_03548_),
    .Q(\e1.alu1.a[25] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _15555_ (.D(_03549_),
    .Q(\e1.alu1.a[26] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _15556_ (.D(_03550_),
    .Q(\e1.alu1.a[27] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _15557_ (.D(_03551_),
    .Q(\e1.alu1.a[28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _15558_ (.D(_03552_),
    .Q(\e1.alu1.a[29] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _15559_ (.D(_03553_),
    .Q(\e1.alu1.a[30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_2 _15560_ (.D(_03554_),
    .Q(\e1.alu1.a[31] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_4 _15561_ (.D(_03555_),
    .Q(\e1.alu1.a1.b[0] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_4 _15562_ (.D(_03556_),
    .Q(\e1.alu1.a1.b[1] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_4 _15563_ (.D(_03557_),
    .Q(\e1.alu1.a1.b[2] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 _15564_ (.D(_03558_),
    .Q(\e1.alu1.a1.b[3] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_4 _15565_ (.D(_03559_),
    .Q(\e1.alu1.a1.b[4] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _15566_ (.D(_03560_),
    .Q(\e1.alu1.a1.b[5] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _15567_ (.D(_03561_),
    .Q(\e1.alu1.a1.b[6] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15568_ (.D(_03562_),
    .Q(\e1.alu1.a1.b[7] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15569_ (.D(_03563_),
    .Q(\e1.alu1.a1.b[8] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15570_ (.D(_03564_),
    .Q(\e1.alu1.a1.b[9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _15571_ (.D(_03565_),
    .Q(\e1.alu1.a1.b[10] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _15572_ (.D(_03566_),
    .Q(\e1.alu1.a1.b[11] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _15573_ (.D(_03567_),
    .Q(\e1.alu1.a1.b[12] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _15574_ (.D(_03568_),
    .Q(\e1.alu1.a1.b[13] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _15575_ (.D(_03569_),
    .Q(\e1.alu1.a1.b[14] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _15576_ (.D(_03570_),
    .Q(\e1.alu1.a1.b[15] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _15577_ (.D(_03571_),
    .Q(\e1.alu1.a1.b[16] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15578_ (.D(_03572_),
    .Q(\e1.alu1.a1.b[17] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 _15579_ (.D(_03573_),
    .Q(\e1.alu1.a1.b[18] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _15580_ (.D(_03574_),
    .Q(\e1.alu1.a1.b[19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _15581_ (.D(_03575_),
    .Q(\e1.alu1.a1.b[20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _15582_ (.D(_03576_),
    .Q(\e1.alu1.a1.b[21] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _15583_ (.D(_03577_),
    .Q(\e1.alu1.a1.b[22] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _15584_ (.D(_03578_),
    .Q(\e1.alu1.a1.b[23] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _15585_ (.D(_03579_),
    .Q(\e1.alu1.a1.b[24] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _15586_ (.D(_03580_),
    .Q(\e1.alu1.a1.b[25] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _15587_ (.D(_03581_),
    .Q(\e1.alu1.a1.b[26] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _15588_ (.D(_03582_),
    .Q(\e1.alu1.a1.b[27] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _15589_ (.D(_03583_),
    .Q(\e1.alu1.a1.b[28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _15590_ (.D(_03584_),
    .Q(\e1.alu1.a1.b[29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _15591_ (.D(_03585_),
    .Q(\e1.alu1.a1.b[30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_2 _15592_ (.D(_03586_),
    .Q(\e1.alu1.a1.b[31] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _15593_ (.D(_03587_),
    .Q(\e1.offset[0] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _15594_ (.D(_03588_),
    .Q(\e1.offset[1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _15595_ (.D(_03589_),
    .Q(\e1.offset[2] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _15596_ (.D(_03590_),
    .Q(\e1.offset[3] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _15597_ (.D(_03591_),
    .Q(\e1.offset[4] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 _15598_ (.D(_03592_),
    .Q(\e1.offset[5] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _15599_ (.D(_03593_),
    .Q(\e1.offset[6] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _15600_ (.D(_03594_),
    .Q(\e1.offset[7] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _15601_ (.D(_03595_),
    .Q(\e1.offset[8] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _15602_ (.D(_03596_),
    .Q(\e1.offset[9] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _15603_ (.D(_03597_),
    .Q(\e1.offset[10] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _15604_ (.D(_03598_),
    .Q(\e1.offset[11] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _15605_ (.D(_03599_),
    .Q(pc[0]),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 _15606_ (.D(_03600_),
    .Q(pc[1]),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _15607_ (.D(_03601_),
    .Q(pc[2]),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _15608_ (.D(_03602_),
    .Q(pc[3]),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _15609_ (.D(_03603_),
    .Q(pc[4]),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _15610_ (.D(_03604_),
    .Q(pc[5]),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _15611_ (.D(_03605_),
    .Q(pc[6]),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_4 _15612_ (.D(_03606_),
    .Q(pc[7]),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_2 _15613_ (.D(_03607_),
    .Q(pc[8]),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _15614_ (.D(_03608_),
    .Q(pc[9]),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_4 _15615_ (.D(_03609_),
    .Q(pc[10]),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _15616_ (.D(_03610_),
    .Q(pc[11]),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _15617_ (.D(_03611_),
    .Q(pc[12]),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _15618_ (.D(_03612_),
    .Q(pc[13]),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _15619_ (.D(_03613_),
    .Q(pc[14]),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 _15620_ (.D(_03614_),
    .Q(pc[15]),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 _15621_ (.D(_03615_),
    .Q(pc[16]),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_4 _15622_ (.D(_03616_),
    .Q(pc[17]),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _15623_ (.D(_03617_),
    .Q(pc[18]),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _15624_ (.D(_03618_),
    .Q(pc[19]),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _15625_ (.D(_03619_),
    .Q(pc[20]),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 _15626_ (.D(_03620_),
    .Q(pc[21]),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_4 _15627_ (.D(_03621_),
    .Q(pc[22]),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _15628_ (.D(_03622_),
    .Q(pc[23]),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _15629_ (.D(_03623_),
    .Q(pc[24]),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _15630_ (.D(_03624_),
    .Q(pc[25]),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_4 _15631_ (.D(_03625_),
    .Q(pc[26]),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_4 _15632_ (.D(_03626_),
    .Q(pc[27]),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _15633_ (.D(_03627_),
    .Q(pc[28]),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _15634_ (.D(_03628_),
    .Q(pc[29]),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 _15635_ (.D(_03629_),
    .Q(pc[30]),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 _15636_ (.D(_03630_),
    .Q(pc[31]),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 _15637_ (.D(_03631_),
    .Q(\next_pc[2] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _15638_ (.D(_03632_),
    .Q(\next_pc[3] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _15639_ (.D(_03633_),
    .Q(\next_pc[4] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _15640_ (.D(_03634_),
    .Q(\next_pc[5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _15641_ (.D(_03635_),
    .Q(\next_pc[6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _15642_ (.D(_03636_),
    .Q(\next_pc[7] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _15643_ (.D(_03637_),
    .Q(\next_pc[8] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _15644_ (.D(_03638_),
    .Q(\next_pc[9] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _15645_ (.D(_03639_),
    .Q(\next_pc[10] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _15646_ (.D(_03640_),
    .Q(\next_pc[11] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _15647_ (.D(_03641_),
    .Q(\next_pc[12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _15648_ (.D(_03642_),
    .Q(\next_pc[13] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _15649_ (.D(_03643_),
    .Q(\next_pc[14] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _15650_ (.D(_03644_),
    .Q(\next_pc[15] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _15651_ (.D(_03645_),
    .Q(\next_pc[16] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _15652_ (.D(_03646_),
    .Q(\next_pc[17] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _15653_ (.D(_03647_),
    .Q(\next_pc[18] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _15654_ (.D(_03648_),
    .Q(\next_pc[19] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _15655_ (.D(_03649_),
    .Q(\next_pc[20] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _15656_ (.D(_03650_),
    .Q(\next_pc[21] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _15657_ (.D(_03651_),
    .Q(\next_pc[22] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _15658_ (.D(_03652_),
    .Q(\next_pc[23] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _15659_ (.D(_03653_),
    .Q(\next_pc[24] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 _15660_ (.D(_03654_),
    .Q(\next_pc[25] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 _15661_ (.D(_03655_),
    .Q(\next_pc[26] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 _15662_ (.D(_03656_),
    .Q(\next_pc[27] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 _15663_ (.D(_03657_),
    .Q(\next_pc[28] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 _15664_ (.D(_03658_),
    .Q(\next_pc[29] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _15665_ (.D(_03659_),
    .Q(\next_pc[30] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _15666_ (.D(_03660_),
    .Q(\next_pc[31] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 _15667_ (.D(_03661_),
    .Q(MEM_X_BRANCH_TAKEN),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _15668_ (.D(_03662_),
    .Q(\next_pc[0] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 _15669_ (.D(_03663_),
    .Q(\next_pc[1] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dlxtn_1 _15670_ (.D(_00000_),
    .Q(\c1.dep_place[2] ),
    .GATE_N(_00003_));
 sky130_fd_sc_hd__dlxtn_1 _15671_ (.D(_00000_),
    .Q(\c1.dep_place[1] ),
    .GATE_N(_00002_));
 sky130_fd_sc_hd__dlxtn_1 _15672_ (.D(_00000_),
    .Q(\c1.dep_place[0] ),
    .GATE_N(_00001_));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2569 ();
 sky130_fd_sc_hd__buf_8 repeater1 (.A(_00020_),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_16 repeater2 (.A(\DEP_PLACE[2] ),
    .X(net2));
 sky130_fd_sc_hd__buf_8 repeater3 (.A(\d1.addr[11] ),
    .X(net3));
 sky130_fd_sc_hd__buf_8 repeater4 (.A(net5),
    .X(net4));
 sky130_fd_sc_hd__buf_6 repeater5 (.A(_00420_),
    .X(net5));
 sky130_fd_sc_hd__buf_8 repeater6 (.A(net7),
    .X(net6));
 sky130_fd_sc_hd__buf_8 repeater7 (.A(ren),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_16 repeater8 (.A(\e1.alu1.a1.b[3] ),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_16 repeater9 (.A(\e1.alu1.a1.b[2] ),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_16 repeater10 (.A(\e1.alu1.a1.b[1] ),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_16 repeater11 (.A(\e1.alu1.a1.b[0] ),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_16 repeater12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_16 repeater13 (.A(\c1.instruction1[18] ),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_16 repeater14 (.A(\c1.instruction1[17] ),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_16 repeater15 (.A(\c1.instruction1[17] ),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_16 repeater16 (.A(net21),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_16 repeater17 (.A(net21),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_16 repeater18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_16 repeater19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_16 repeater20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_16 repeater21 (.A(\c1.instruction1[16] ),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_16 repeater22 (.A(net24),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_16 repeater23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_12 repeater24 (.A(net30),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_16 repeater25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_16 repeater26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_16 repeater27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_16 repeater28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_12 repeater29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_16 repeater30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_16 repeater31 (.A(\c1.instruction1[15] ),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_16 repeater32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_16 repeater33 (.A(\c1.instruction1[23] ),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_16 repeater34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_16 repeater35 (.A(\c1.instruction1[22] ),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_16 repeater36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_16 repeater37 (.A(net40),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_16 repeater38 (.A(net40),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_16 repeater39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_16 repeater40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_16 repeater41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_16 repeater42 (.A(\c1.instruction1[21] ),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_16 repeater43 (.A(net52),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_16 repeater44 (.A(net46),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_16 repeater45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_12 repeater46 (.A(net49),
    .X(net46));
 sky130_fd_sc_hd__buf_12 repeater47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_16 repeater48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_16 repeater49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_16 repeater50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_16 repeater51 (.A(\c1.instruction1[20] ),
    .X(net51));
 sky130_fd_sc_hd__buf_12 repeater52 (.A(\c1.instruction1[20] ),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_16 repeater53 (.A(\c1.instruction1[24] ),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_16 repeater54 (.A(\c1.instruction1[19] ),
    .X(net54));
 sky130_fd_sc_hd__inv_2 _07523__1 (.A(clknet_leaf_8_clk),
    .Y(net55));
 sky130_fd_sc_hd__inv_2 _07523__2 (.A(clknet_leaf_8_clk),
    .Y(net56));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_1_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_opt_3_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_opt_4_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_opt_5_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_1_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_opt_11_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_3_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_3_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_opt_6_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_2_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_1_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_1_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_opt_7_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_opt_8_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_2_0_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_opt_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_clk (.A(clknet_2_0_0_clk),
    .X(clknet_opt_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_clk (.A(clknet_2_1_0_clk),
    .X(clknet_opt_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_clk (.A(clknet_2_1_0_clk),
    .X(clknet_opt_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_clk (.A(clknet_2_1_0_clk),
    .X(clknet_opt_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_clk (.A(clknet_2_1_0_clk),
    .X(clknet_opt_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_clk (.A(clknet_2_1_0_clk),
    .X(clknet_opt_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_7_clk (.A(clknet_2_1_0_clk),
    .X(clknet_opt_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_8_clk (.A(clknet_2_1_0_clk),
    .X(clknet_opt_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_9_clk (.A(clknet_2_3_0_clk),
    .X(clknet_opt_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_10_clk (.A(clknet_2_3_0_clk),
    .X(clknet_opt_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_11_clk (.A(clknet_2_3_0_clk),
    .X(clknet_opt_11_clk));
endmodule
